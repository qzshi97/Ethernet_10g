// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:28:47 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SZYzgN/QfbFuS/65i2sFIpXezrmOmtQ4Dly/iCNwAOARcfqUvhQ0hNmT5+ycydBO
FZeMy3imjdN+oU27FRhVBDT7iczKuv5eGeDm8Bq66xzXfFqteVvzw1zBt3EYzLBv
9cicM8QdWrqVdz3NRW2Ewm6yarjU6HS3Ktmr3q7uZDA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34720)
nfxlOKc6Q0a/YPW6DaOsftWMFaDpMnUyd70Ow1FwlOHq7nMGvJVX96gX7/oVZsKc
Rpm7kLMSvCUYUVrL+XQUdDUzxf0pNI5Xsprn4hj3FCv1XxDksAxxCx7JtGcVorUh
Po8I3iOr+PlxDAkMuoK9iCK31at6COTZv4j99Amw2CqIJ9tOp11rFJkhpXwrthHw
SuvpbtTPQa6EG5ogXzOFqRLXR4tjlPCbunMoHYnK1opbp2f3ln06BeOukAhsUAnL
hXh3xUK+8+BvLDt0r3lHzPjVRQOMnPGI5HZkxIhjEkkoTQecdxOWIIudARqJqcmx
XusbkJHenjpKA5AX1DdY3OUCQI8T8JOyoNuTxVadiZdBs/ERt437Qd6E/elKcgOP
3ByxZKJvujtpa1t78RQ580iruCDJtURKS7OG1uudBDATtXdj5r3esvya20VowpGg
3dh1QTIZ/YL+puivHiC4XQR6sI6o8p7iRiEusJBMblv+z8XgVkSvBeSdYQT6hdjx
ehrpY9quiTbRWtN54iig3B7TdCA5AhzIT76RgsQb5lnSzgCLHXBZzuvvr53v4r1r
VCbImk/YBHbIkxZjsmKO5gaMhU/d6t+1RZmhRRREOUxssPPAssbIoFc73ZdDuTDC
t9XUzHQ8Tf68G6Ly+tJWTbd5va35+0q2BRev0T42pgUuBEv8+a60ktLrQxtX+o+K
AZnDmNLgjsPVPrbBelEhUeKgHNNgdUReTnBBJL0NCju+ylk9kxUuDz+aRCVUJGRK
y3VVnHQv7948jN/UqYeIWbBQRo7JYgOyuQ2cs+oQhV19kcGo1LzigQmk8Hn1cb/4
as5jqFD8H+CLlXJvQbNX4IpSChEK3uhIkoJ0PvzaxPjQSU3ScMIL73KrV20xG5wI
ji/e02YPlnO2nElx2gn7GNLMpnOAh8/4w4CAe9JCfGeQXEZbO4FoEDpcpP4BXh3o
I0lnvT70I24Ll1FGzYbnYDtXal7CEf0PlSf26w/L1/KUzPy3ykOe2/3sexF5+u7G
GPFNOKb05dpqIJhqoNlrWSyPxahoz3BovPa924KSVbNjz2XXAmQUn+K33D5z/aYH
DhGsrZf22hxcScx85sfYpJOmKzWLGvce8r2Yy9jgQNPcDSGt83H8dQmqqgMIx3hD
S8yjTWpkSPtkiJMuqeNMUmhPePQe+1nU1CAGL7s7NXVXlRbB0KnI6OFyjmVM2L6L
Nrkl+k8TbtHIyrk/8XIlBj+KS20LqDYzaGSS+2Lp64oHCbx+QzG9W7L9lMe+SUvQ
3PM3h5jlC0ucugB5guu8Htd3P0v2LIeMfS7OLkobEfK1vR1P9j1ICdGVgudAof3V
dSxnxBhz+1b+llSH5tyyf70xXto2fnLokEq/b8UX+b+kbHD2TlyXY4RraXI4yi5K
VqHHtremB5NrlQTIv+w1UDBRlrx0CUUFna9GqXO7x3DbBeLL6SJe8WcsER717J41
rN8mUKy2747JrNEM0lprrb0aE1RjBHh7+o1RcfIZGrU3Pff25oakdTPZYiHhXE2J
0uNDqkZjRPZ7vBBzhZzjYYqfxu1dJBh0OAClrvUV5/myhHhuwKYbGXX1bL2R6Ks5
FkMpSKE024TzsbYRu9303BdPPC/btRR7rWnwd7UD1Nz2oUWOACn03STAT/Y/T/e4
Ljybo8u1BiFWyNVnXdq6TpVT3YFQs4KEIpg1WDSStP+0YzOq8Qs13QYMbyu2PYDy
yzRAoDMVEizNvzu1jNtB7osJ0KzBgmbAn2fI2+VlYg5ZQ/5Iu1IoADObqtD00QvR
tykVa06/0T5VtXVe7osEWNvRje1XdXzHR+4t0NB3NwId7acSjG/dFZQQ95Sqisuv
j0Ii1SE+vN7ySKf5F7gnryVL+HgRlcvZRj4U2MrTLvqfDDONaaUJCuAlzpNPJt+/
7w6Mg2InAz9NhrBQ7KadrliOPuKjBsQt6NwtrKBfF9/JURBItAFpoDCgvj6bUKm4
NeHKU3POm8kPiIObq/6IuWBEpqq/cd6RpGAAmTZyQzrVo0VwhSX+N1Oz5WhLGfQK
UY/NI2FQxwyDYKycN3gkTFqvidPSm6r9Lpw+/nAsA22L9AkCQCYyhWRdJBJDerQz
FuyGkHfu+C1lfkmrdkyE/8R9AbFN4Pbb/Oga8wgQd5SPWhzndfVaZgct3G9wK51T
dqTT/+AFJxCOTGLv2l72PRAhs/r05bxQsPj0Usfx6JJH2mZn5QdGZ/S3K9jbXCCZ
fcETR1l7wuRacxDzWGjTCxRa1pTzzuRxEV7PAw+xbFmGAvYgxZ8Ag7MTWaAlseRv
LNo32ZtXokqJ3ZrxluRALh5qDYvYavimEYnrSVbpG0dAsrV6tRYtQsgoj6wyC6zv
EpElhl+5DzsKtYvZJYL7rjW8sklhEe94NS1Qu/yCZ0LfOm9XnIfEE9tFXlEjZODK
HRLVi5YTyjGFV7MmvLKeR2nLiPA1H3xbDfHZXE3BuDXsnhoGgHej5wD/KKA3SLzE
c549nouqpZn9yhtzlubWAgxLCYpkbtw4Q7N7O3lpu17rp2N0Xj2vecHZcpvVw0/J
yoFR9CoimUlZlelJcC7rKw1BUnzecXiUj+3lZaOcz9l74wGwVG2jbQag81tWhrOv
6lRJ0yR+dxia2KsmeXzfVZQrtCTq0QqpfvHxMN/LHtGDj/Ru51cPgcCiA3naKb4K
JEypojBE4HeFXHhElw/QXFwmCTs65S+u3BI5ROb9vC6oBfg0XxdLMrD6J6EG/KYS
wBtnd+0NGPsac/ullPFH8FUGbjQRX5+EqHqk6c8Y5SS5PXui9keeidRXTelhF4oh
db8yaZ2Bs87S9LAmkFFlNYlZ9FA/AJN5YCLYdh0GzMkCZsf/CLkDQTJWMbOKE8VH
3mFD0r/Sb88v7WzXs4yWOg5S7XViGxpBl0MMPL9x5vLe/lnH/68lsfbkco362oj/
t5YogK6nuC6UBw3teqw57SISVWTjFsnvnPhVznGRGDohy0TcnOajE7q1l3LRNK5A
9fohvjaysywytJSimBxGryOjmMaqIxv5In2Y2rkh7qR1vKuQB3ZRjqFzfdluXdbe
MqCPFDxQePE/ovGonYnvi7FMMtqe7X3W4UXPqTxanCsiqVo2nzxF96M3C2I9hKI7
iwZf+0Lv3RM/Omo9Fbme8cdv0q62OXTIpk9pEKIlTzEzcarlVqnMU4oO5sYIctk4
9ian8nq1AhynYskyRBWLKX0um52HL4wbiqvHTI84RjYXXcv9m3oFq+f8yDMeIntn
mRAD+oJAVwPmzTeSL7DjQko9IA3eOMuAGWqlbKeggKdvZpXJoA6tlz+i1O+t+R0u
gELyVrFGzpTN3GTBoEUqrxtQKnLmqrPb86Ix+uL4pKxXOz1XOijNzhG4L33xG79v
0ij/bP+dwyyDOC13e/S+WExj7JRlKjTAI7gtA3lAZJu4CR7ydUIvH3G5scy6jg69
HMOcuFFN+Q1JkmPOj7e7sM2FCoJWXIi2o/Ec1rL0iksBkd48HeApRIIF35VfF+Wo
+PszSYJoESjovw2bOtGrJ90eGrDRczLbpgamN2V6TScxT7lmS41MRUQi3m0B4dUI
xpgLVbiJ/n+aWHtCSKgih8fHxahhX/4o0yt7QEL4oMG4iU0XJKGKGPV1nrQXx8wh
FBf5ya2GrL6B9xPBvzznQ9fa1Y1nNSPTb/UAq95eKDpEwfpjLG8HwHe9kArTDs3T
w5APQsRtMD8HBmLV8Wzlb5NGGxBxgvalha8XIIy00Nm56aY4K+nh0MQoqiBM0m73
p4EWDJ4yHd/Tc/tYAzO74jIc1QYuP6Hj0cS3K1d1d9bnHf2n1Ouy9bjh/UTDsx9Z
XrFGjwnjMRd6CzdI5CmQTDR549HeFUGtoALcGQpC2QRi6jFpzFh/kb7gaGk86p3Y
0vmsHrL+jH34C1bGCMzWGuK8T1t1XHHdQ58D6JZ3dvMqjDpn1Aa/ktp4E02k5xYC
0dkqZ9oF3pFWwU0q2e/IdXXQzXnA4hu2z9bkR4hATS1UZqlZ3JeE2kSd9LwvHZP7
VyJXtYaDGUrNsZTIPywuR/J0QVTjwlsQNVSkLOsGKZCqNsiPqk4PJDvdN1rMPkFZ
OUlf0rNXMJ1RaR//7Trbv4bgaB2qSkitOTtT/O+Y6vzae/3EHEVWPYUUaj2PWAmV
dAY5a54KLcnYV4zKqVYxfEhOrTPVSltt07JB/o/ACf5D3plT984p3UP7IlM8hDkc
OsFHxSNqpCTHHLdGNHR3neGAEZ1q96izp7z3QIJbvmQwjDLRNhaAy6ImgTT8cW4J
cfQ3btbflJHFYeGjJWEWkhr97LEae/yNLtlOgihMSh8cN5rFhz2fbodMWcYORQIi
Xv5T+wEZMIhQVAdb+sSuUWxhtdB8JAZT7QJiHkBdctNPXuiTZp4ktsfzHoE2AZOs
JO1LyMU7pAwUz5SMAXtfW+B+j3m274fUQzATUVO5FSXvHJAHUE9t+yL4kO2CzG69
uiU2HiBF0RHoGGDpzm1rWw3GgWQEU/QKhnm5IieqUYFkZAZRz0xcBet7zWWquX+4
j7hXj15VrUU+qbJutvaDKEJ/M1DcRN8ywIA4QFh6SxRDX1Rg7VjONGH6hLsNpxwP
uu6FVtAsbcR0F3TO1HG1FQZFz7TprCn5cNhmSdq+jnIku06MXWgkoDqgmZt6WSz1
nn1wPD1rjk7xqzrKpFqFjzNgqhT6Diyok432ujCue5C+bqk252/EAaeWgPdbm1wY
O2RDL3QatlfIuY6uTcYYohbQpz3dIVCXkGQuqFFcbTWksLYRyYpI1d/BPvFMle8+
x41Ynt+C5qMFMqAu+t0SaZHXaD0Ujsj5oqJXvRMPHFeZCDPlQPWir43VL4u8QEAF
Uy2ODrfQBM0bCMv4X8+gXGeDEyfYS6vVWnMjblU2bcm/cw+CJ5SsRDHyQ/TKH9CV
6E3NVPd8X1No0iWw6riqiyBWAmW03IMHBYimZnFdD+gJgXv48edwn+estCSVnf/t
nmwHDr8a0QWZieTuXg7S0XWvXmtT6q9PcBCxct3t5/9ti1rKncxe8lFLeE3Q4mmf
qSXyq5WRw6KDHnGs6+QVWdiPCNyuKVyoj04bCiEGJrmUGsPmOOT8RH/f8B00Ff1N
rJ+vdyzcEwrNS5ea3IKQ5n4YW4uZchfxm+E/Ms2pQ4NPcBdvAe2TjAbtxjd5ASMN
ZdgOeWl5Lo1SDqnIGPsECSzDt1SIAo4/pN1qJUHwVpWLAS9k3CvN8ujM+7Id2QHy
Q/fZbV2dpsp930yHahp7148J8Bt1Kl0rmWnNnxPCyhbBJ7lrkVAeBjqdpp8YqSfv
y636XSCeB5usjAMcmnC1DywMo8Xg42m6VG9C+wK0I6BX/+7YQkuI17NkDYtd8nr2
usGRSXhTZ8/sgk6m6/CfKo6J/hHF39KJNMJcR3kA14ufDk/SazrQDIb6KDhM1iTs
MSET2annTkxU4bE4UNrBS9pGp055XCUeJS6kSBvN7WOspI/G6YXsjfzL1MtMacOj
Kdl8+e8RvGYfPP7pBelRuzzyIrbBx03AaWT2THkSEIURyJAHCa1Sbfjdv0oc6CQp
nwBSUgecD5FpYbZRCMZ+PTOz0/hDqnnZH2vUXR9jXZyjqdQUKDvlCz0ogreXa4pn
Hd7k7ir/e/KLMiVdXGgT1YnEcApu5Div+qLCBi/+BZ+ZixHM+QnQ2KUNvXwzffeG
X9Rp//58EywWIAeg07923AFQSEK8G/W4grphYXZybYqfyHn7BUNtIOovcQ7Yb75D
anEPV41xLyJjSuFsiZ9rVltTq3cJ6hFO3ytH76aAf6inOYpcBcWC0k0OMN9QQy7z
Bnl068PoU7YuXKEOicz7YnXrrjurnQ6Dkk68SLIXT16hXy4HRHH3bVydKvOLiZUl
cV5VRdW59xPIO3Bo/MFhDbkm/4xPjgvjs6H8TUtehYcRbKTfUmB4DUYoXl8vSCme
intAOjtf+yadNFtiWykWR6ijo1qc7s8UdVaeeItX8A5YwwKgXOSmpwRkZl2S6uji
o80f72JyV8BCT0XGXhLGY8d6d60Hjy8+PMnAPeNpFkNtODT8XyUXLCvoqZNID932
b+dnGKPYe0eFbie+YhNSr3svqKnGijZb/J5ax4IWS+lggBssTxSzBz6ceuQ+yrtC
3e0uFTXHdSojKVkehpTl+GGLOSw8ikYM1PLfq/1PtoIMpLQZ8HdJzOkFuIoIP8Kp
euHc7rqHvlk52Ga6tbRz5x2WewNM03GxdwahZTC/lFA0mfqyN4K5MtPABzOS2OnW
iIVH6CWS5j99Xcv9op7f5qmDbgxlFlPz+1WbZPFW4GBIMYGV37dlVkkS8LKvhh14
syt0VJtWgkgjY0W89TU5K6QtvGNtFWHC5MrD+rkdfv3KSzTCQSMa2ulSyaCXgZ5m
YElaKEZSV+Ah1Bwbsh9OO5DgCyjdH4GseabjL1Q5ZPUr0RlgnZTNVwDrvOT3MT3v
lLUZ5YdNydUPpcmlF/av07mun8QD1JnlWurj8Ctw06y/NZsVlO0ITNEj1w7H6mrO
gDnzUKkxmzr9VQwizJSenrEEwU+s8MqmsY9GErbnEkZgXWSRemTARej3Ls+Z8vdT
qZZvqmjsnQl1IDBLu71aXnujTgo2xPZTx0/PEtcbm3H3kC0tykhjHUJXMn65qZ3T
KK6QVx4NfqtF0ybv3dyQNpQJI1vNg6TkfB1+uoAFys5grjkd8Suus/hzXJkdkICk
edAEqG/7Jcllm5hcTY0EVjWBc6/lDAxfB+Hm0RiQJz01dz+fLPKRzxsX8iowzWm8
LAGEhNyAuoVEZ9D74Dt02SgbzRwWcWatc5YnSD1FujzT+LYf6ATAISRzD0yQ1vFC
F9xRC4rgIB6Qbj1aZ1ZYOyX/OApKbQMz1/+ku7JnpvuP/3Qxo+iqrsjLvbMPMS8H
Y1uZ5iLiqYNQv/Nsijo6TpS6VZoIjH7O/Ll9Zw6fjTovqHIAdhpGh6UnHcFheZ08
IdMaMmFwBNiQCkQxtvUb9iSfGIEEo+Djfb3vbZKMeGl+cFXolckCx0ZSbEPA2c0Z
B9FA7zOSb1onxywN8Gv95k32etHrzjBqHNt3a4I0QZTmvKNNCH0MrtoXr/j+NxE+
QOHjSzq5UZgzurgsWwB9pKYogOLPXDRqKe2gdozyvG795i7SyJJk8q/nvT3F6QbA
d1jACZjTvWWyKCRC91dSKeFmsCJnnKD6rAtvp4s6j/4Cq13ptD8T5MGs4JpSuCkU
S/oaqaa5XW0L3YTH9qEGMf6QYpwp9eki6JIrfE9Jt0hs2LJ6KLnJ/vQYEKVVw4xK
ACsrSnF9UOFJ7YvAxalogej1pgaOodIJ8+tS3WGz7xkiT3yIo+dC4idOW1bfidSc
Ywx/9gO0Yx0FGFxIOj4PwuzzUFLpnf6IIRTPHA3/wK62d+US5JozFPkDGfTyA0iz
ssUu3CEZ6Z4GYEY54lhU8otRy4qYUk1V46WcOt71TjhIQRHP1fTbl97OEMf+HLTh
ecMLXRufNP3qDVvNV/PjXhEVLb7H3VJ2ap06VCNkJ2oBfRSBMkj5C5JzUVMq3EgA
rUJWKa1ZEj5mx5zkcjQReA0fpT/dTZDB9ytf08/qhp5e0+C2bTAzGgBK6mKCbdjV
vAkZq0Rz5E4tIYXfR2IjKSxEOSdTufYQ5HRdw40VtU5gnf6Td8B8XvwG8F3t8qlg
NO9T2X2CQBHn9hoeYJ+hZoPxFFojejHr/g0xtpZsloqVV2/yj6xrzdKxb/OflZzs
f9oqSONwImiyg2R1jeowdhbe+aBS6QRMMiIMUdBEvbMHWc0aCxMoTN+VpBTWntUC
uKLtTKjiFpiUffbxjFXyDNXEDZm0TFSaOoGcOsm0vhtMRm3VGkDHXGvk1A6oYyIB
PXpFxIhOWvN5NE8DQc012uHSn5pBQdmnSZaVf5vur33xvSOs1sxW5/6DebSojkLq
zebW0TEGIPKCx6L6IFg2+hB8/va1WrYFhXZAThMY5ro9pmTlN7mAcSfgRsU947jV
fUZXjZB23CJe3CSL+KaU1uHOAFScmzXCCHKwG3AxAp3XReC6qpYS714aDeo1t8nZ
VK3K039osFFQMaizRMLbrjoQR8sVhCmlluWiDxHikqZox7CLRGrmU+59xG8mV2fv
tPtRp1TVh3Od6gVM/2A3WMx/vn6O8R6igf6SjuMo6CZoSHfJsxAVtyqO/LgmoThD
Zc15L70HjeE0i9auVgrK5xEU0zsq6xFEMLcY2s6Jo7sKuf6DHZFK/mUPS3sXrSEK
VQwd1oOqz2MoLqUUMvwJIX4bJConmxo9daBSfZ1iEhI4Z1fsfumA3QM/bJtQmjNg
ZMXui6jkxELkQMXc+m4TK9ZO9hS6RBpVUMM1nh9s6sJel5aUd9T/6WLv38brHdkB
zODZMSmdd+ROItUTG2JP4jrtDpp/loRZidV+LcPt0G+U+OQa+mQn1hK5EZ4u2d85
5EZgQh6ljIupPEBcs4QIpD5CJj7RIX9TPt1dr0gN78TTE/VLqYGf3p80CP84IAJS
vX0+KmIFDG9aubvNOxtBBWX7lE/NemzV4dahfjoj9rWou5C/HeaZKn3C+3sKGzWz
ANOIOhh82x20cMwt09tPb/ZKz7/gkx267HQ38ydvHFUBtYKAXnD5UrUG9w49lMNI
rQGdaZkgXphtBwA6E9yLnv2mtrp/3hjLcNETP75Fgc9MdlYiegAJyOArjBTvks6/
OhpdVYj1F2aY77G3rUlSi49plBfE1NzJtzDdrD+lZJiubbjQoUJeZtDUkBV3yd9A
LNdUSn9wdWUXoqlNhbqsgjdxkLMMz1Gx356FP5i2pT30Al4CFlwl+P8uB3XDBSJ6
y0cBcgPNHUjYGz+xSm8kcnVXL16ZFuS/Q4LqTW6Zonga40/Roa3K7R5ByYOhFmB2
Lo3hXoI07HQHTlgJ/HYeqC4V3Pr1Lj8lOFe2hiNioY/ckLrNXRzNSKTnVmvbuhDS
meCEcZL00zXXxhK6XyO6VoHI5hw/PxlgrSOlhoyLSSzx4cawK+u/5xB7hyHlfX2s
/w9kqzaJEBxqyGi25U4FGsHB7tWGDBl5XGiNGxV9/thhh98SrNmAvMYku7TfDJkN
ai3vdYpYJILQDvj4U/jcchFrjBzrd5dMR6KqUKvlLf3tXsmz5AuwizFhBW5brtHe
ZO3A3gyWG9RxEC0bLMnhRcYNPLMSUN1v9MmNrfhLPrvyNuItwiiBBWRd5hBIwBk8
qhnuIjNd/yslhXAQD+GTO3TBblEU/7BMu2j8uqGuFpci2o6tErWj7Bv/zNJZYhei
iO3xnXxC1BisdhBNX8TR1RofueW8cVVmkvLhnTsZrKuXS5zrmznq0ZBxicnPy8hS
m7YzVNZ0YuNUgdqH+a9OQT5lgTF0nGeYVpS1ov9GTlUs8J1mvRPYmTP8ISjvkWiV
uXfyVR6WXJEeVPv0BpuNkvn+nHmfQTx9iglUTIQFGA/Sr2XtnKadom6CHD7qmQhe
zNPx4Pl9wynjn9S0H2Jr0XxFCKUND4tTqCF9NsR6KyxwyxWMdAV7N7Z9UdSa6L7c
bQ84GVuBFeZG5935nEBhsOmig0MmbZOesCdHQ8b2DC2ktMrtzRbivNpOyJfbIuIm
WmaVxKxEFpiDhR1VoS5xTPomMdpvhwWK8cxjkpWc70AzXtznLU2K86Xucmnh78Kl
E4TXBHvcAfPLIqxG6Cl2mZ539VSHohLYmrrWzq+rV96Srcyj3TuoV6BHHXj/vMr6
6zymC6IhWbaxdyHycjPIMY31EGlghC7rusYlTRMlQw6h7ONCbGtMI67UHoS0VRsE
2HbMPpP9OEOJ9KrHjEvMfQeWePe9piyhj/CLHn+GN2ho6lTSYbyN4pusimryZUmO
/ALPODOI2ymd5nj53X85WF2nsjXA3FbT9KaapmAuZBvxJ+emCf41aEZ4gQida/Yt
uAMfwtyKkc+kC8jIB7OcTFWLNy5SJmpI17WkAM1NiEoNkTpxXqdEGc2KCQKP8XK8
hGIal2D60LW0MeBXck9MZwu34uMBpID7P0f/zdwHqAtsKfEE1V4P+F4+jPheTb2R
wneVPGO6bm63UEcCh+F1/k4eYl/yiQAArcKrnNgwbZxQUj8aUYvUC+53Cq3LDzBH
YJA7Uerva9disJSJ7ZhCrCyVEWsMJmjQx4DWhVw6Gerj0t4BUkDh44zdoC3MVbfi
s5AD6yOoLg+iFzLjnvnK2WU57pEZHKjqzoiM8vIM0BaCnRvE3H+dcRfnoWHhxlp2
Ak1whLsccDUDOhi6ygSTr7zgaty+rXOThoBRV9Vd11/gYmqgwOupUAr2mhKVhWkF
09WxIbYCEc1apd1rGphMPeEBiqeK3z4UkIpdgU99o4bqB8D0SVbHHNicTRmZ8eYt
RVK35BNhrqfeKBYn1frcTXZTf0K7AcTgfO407ZOgMvm5JJyrDQFPxOBTphBfJWLH
rcWuc9m1nUnOQJUDmzYSlUzjqFQp/v8fCP3XUfez6C5Ja49tuUbE+RdxPpNi4/gx
C4L8QDeJ7NX/q+Bkd6aYczi6+sd7pFSnwKgPJyOM9GLFFwITzk+DjTxi06wjcXuy
PFHnxVrP33sqhgJtObt6ShkIHdWJ2Blg/EKRV7qNCcQZz71+qEdB0ULrCAq8mtNy
7GeuEnYOyTZe8tXYayxoYtDmoy4apKW1aEtg4Pq/CbJMb/nV4gtigulnBVzjUa8q
fcLzbhCU6GS20yIjseKaWPIpDGBgKOUxwbDFOyP39PKbesLFMSV1zvJAQ/xAh5KB
MhmmganWqn7/TfHKXTG2fjPiY4l5ktHMfF9qQBYzQTjffbik2H03GMBYHp5pNK5Y
2Vt5HElZ92tE73OEnhcnNaLJaPwCEjljqg/GCeRarze0TlOq+teLRI59HECyzlPW
AvJmOCsm4JZqnXosuWvjMDHcyju88DRCwkwGhO6CVy1B5HJWlDNCsVlKhdPNicsf
yijSM/XtFOZl++o8e9jqldqznQAyyiLSu6GtH+A6zQnwPOI+OYuMNLPHc+9LcQ58
IpYgTOSEYRTE3oO9fouo+xzBsKDG4h/lpcN5RUp2jiHa1i8RlbgDAZAr1XtdkrzT
gYP430++oGKkt/CO0pK+DMOZBhs0i+Mt6kFsb8tZ07+jVZFEfQov9WLRfjHHna+8
XUxrURN2UODz4G1f1rYT/xo6sjRfrIqyAmqYbyB2MZhjuDcz5Nt4Ln4gcaqal3kP
4OM6WWt3p96ZTu4jtAQF4wRkd95rqbCQRwdvSTnlQMs1JYyIhIV651KymihI4Zvq
HqA/mcK4QAG3i/B38CY7DRwK/Dcaazut8sOXDpBD18j70SiMYNX7A9CeqlBd+a2O
m5ikQQgbl/dZz/wNjkNOZWP4uNh7x/tOZnebcuujDAW+RcKxZ9Ecw8Ud4OMhmuYr
d3BH7ZP8CxQ08LenGw+ClvRMhRWs32EaKmcbCADD7TAiqRQxouG99G3IkFaxO2dF
d6UQp/+35pU+kCElKUP0zpE4A8qZ+Q94+sYc/1rb01ocPhx2PzQDf5ZVi95zq3Ci
GTpFL6kQyWLyEwd4SU4pQyMpGoEwfm2uZgGrJvz1+09HxbhWk4GOaVr/0eMGW12A
7px35VnPP2RD5edvwNQI5aJeg5YH83ab+40jw1n4dKkrR18RzW55fkHdwK3/UROR
fO+tMProy2VvUsJAosDSYnicZZWSSjOb1SVcqffZ+vXbjhndXJcreikKSXRrhg5c
osnXwItIppe78RTqA8+ErOlkaUdUfHKfirmMoS6hW0T6/W88r7HfumkHkHfUctiD
xQvsgJmhT7dYYQldscERoL0hlAChIBHnPTtg1Ptd7bGlLJVrlPhvJ5k5fvT3qBWM
+JOTjOURoQCP3Ci+o9d92z1p01Op9Ui7o/KszBo9nohhIjZkVSaV0o733W4UHCW+
hFI0bBzXtOTYkaV2rnVqOfa53SmuUKM1BNSqBUYa7XV21c0nHE4ACou1SMZ9FUkd
toVmGKUMGdL4+VYRykNiLdLnqv2fpWUIn7UFsuvcIKKHJt+AP0SY/LbGdpogVt+j
aQQNYw885Rkh550zkWJ93cqREJHLlSB5tKenNp056AMncn8Hl2On3IcrNJr2tQc4
Derq7KqTKi5e58NIDi/4ogRl9qj4UFDzgfgGZ+YxlB/llp8t29NCsWSm+ZUVeluN
O0Y1f3RIj8f+/K9Ow2s6/F7m56S5/dciin/qsxeQj5Nsg1tKy19Qc7AmuctYdXPh
6Sq0QUpmEXyQTZTkl1k1Wp4Zma0IsF+YI/jQcWD7J+jwhVTSKJ10q70D7DRxXtYO
QXvQF4Wtc59YNear33oiFzDDVt9z1Ac+PbNuTvWDTGj2VFxutLBnBYb+tEEEWAiK
Gx7UrgGdcfvXgtnWHMMaoGy3+bZsCZpa9FPQncIMhK1zqx2XYWEBzMfr0RjF8ATu
pmIB3DCUceZpE0yNzdvEOl8lzgkh4HSBjCn0rxs9Hb97wFW7hLIArVt56aV+19he
eCZJx1S9jyakrFqfCN3VJVYQDpQTDipxKhFnje4d/Bc6aER3LUnzgYMznmwU19DN
u4EvWiuCL/5FcAQEdK49z5PXnZzu4ExRwQFb1K2lrIeyRORrrX4Z5l3atwyweaJJ
ruxF+UVCDCWlNv5/omxOJf7APYP3mZygV2jNBVcFj0uFQhCCu4jRMuuZoALYL1fw
lsl02FMKAoBA0CFztONqKdrR5rb1n72iFVXqzl2xkRF4EhcjScfP6uuNEF881Z0Q
BOjInCzQYFk4JS/bi/Xu37MDPMww/A/MOeWO3tRDbqze8n16YdaaCHFxQ+ER9Mf+
WOdhLCUXDu5tHyynC4RAaoZiBHuNVvAYiZlRjD8/j8uTqPdV/Uw+DePMmUe/45Kn
wRsQingGi6OWJ98gt1Smqh0OJExu//N9bhASvwvyGAutY/6eeHSSCJp3D3rdbbvw
vSIHe8eC+5FZU4a94pVE1yx/QPzYSoQMCQfwAhd8CChIM3ytwLtTJki5taLMbff7
BcOSr41Th5f7Z+fKdbkz3jixFQSYbMVLGJfUSTtT4H0Kk9+gYYtAfCbml/GPbBDe
Xg1VgJhuROZKUsP5vm7KJbRPiO5q5+G3m1YCXd98zV188vJkNeyFE+O8sjOtqTMr
7ttluHx38eFHJw7ZZa4mrTn/LritKQ8EbPP/6tLFGem3BTc1VcG/Q7YGmXfFshKc
NCWNos55Q5UCQcbdchUMFFkFaBjfKN55Uw8fha3DMxmg14+HFIwQefJ8kfuS/nwn
Km/QuLUy77UkXB+/hEMcuhklPYxlrfCH9vUDTshUItTR+08dSY9e2LAJJ/F1oDQE
r1kZS1gHvn+Ln6FZWNTBnAz9rDZGglwL01XBioYOGtWaHQeFMH1VHguvb4y3HMNL
78YeAuW3BnWoANIYTNVnrgKrC0Y+BK7d+Hn4ZCjRohpkL4A4IeOHmb7Tkbhgc6rw
ljKAdBv3iBf2GBgfVhvGDkCZUmqfuoVS6kSWooV9jOHMrTv6tBzodzKEoi7uzMz0
/9jEZebqHwkkXsBayuZ08nMeN7qOqhD6B7eorn7ESXCWp6dTPiN0rq9H8feIRky1
kIxnWpXCAUjVyfglxSt8vKsCdQGm1oqA14t/AtbOvk62cUYmf9Y4HTXIcze3pZ8u
MYBMno8jaTYJhjPgRjE7n75dmQXgN2AEJ19+hG4YTSY2AT+oI1X+QKC/Kr8Ieldf
1ywK2upzbudHmhqg7iA20DRigrx7tKhUhecKE3fFkfJHgJMmXqezkPbOk3F8siS8
gaXjJE1nFyviUOCAoH7/pljp8s1I2Cb2jKgKfmp94Km4g4XjzAnOduLFH9Asgnmb
hEFIvkoMwjUyd8A+cB/CfrKw0re+clvqgsNK9EBMqECZV8MWd/SWoNdva1f0dZlW
Eeen8iObCLBf6/jiUYwZQ4U5XL2yQIE+XE78+kS8VUMoN6TKqKOpcuWjuY9VkiAI
eZY3+0FeM7Gc47Wm9AQaiycDwtdRm+wuWdFmr18GIuvQvit2oitB3KkwDy7WKQER
9NGL8JLXCnBR3bLDjaugRCHeIdZeLC3F9OyLCSdoC3T23FYvtRIbiadYYogGU05r
cEUuP+5DJcuC5eDoKW0ViNVjun0WUpeNdtnQJ+hI5KgwSr7g0SMAQCrMgf9ri6eL
ZIUY+Q8ADPVq1U9bK5WbFel/NoXGt5q13uGKs7hCIE00HLGPNsOkVGdoxT+noIWi
CtCuC97o6GwuTCGbDrfrPVXER0N1mgNjKakRIt/h/JAZeq1EYhktsf3kaUO6GOst
gGDAPJTw73wN0VuCK4+aPOtKKu/0l8KskVSNE8G2+7fJLgt88Ewi1bYyUd4LphcB
Mt2mmnGtlPhCHCz9YFgFZA1ZD60yPILE51HzFUi7jmgmptDw951U2j9wvioKo1rH
H3xmko9cvelEyoE7aUqKDRI7JaxAwTeCcXnbmhpm/c4h/GEAxCI5o7LHyw6myFp5
xiMOIy0NklYT3wsB2MjzZVE4imowwq5Cq+YRF0sGTsBD0AKff67ebFOnkUu4hKUp
urf7QeBFcs3OdZOlRavpsCLAARLkDj4ierQtH0EBSIOxYw92IqjqeeyCNT8cmpPj
QE0uo8IJXKbbyLMwTkSRZyyuHzWrOXJbDgjenesuGsek4YqKMu6oyuMcMJ5BFG16
69qDTt4o1kpTZYVdgDXjiDKpz2ceHvN9Xae51tjqjMGRo7bXH2RBGiygAzwj+XmB
Ee8aeCXmSgz8O2vrFFxbZNKKkDzWreVMx3+u7FCcAQCjKz7zmFI7WobXNZueqTU6
1LqOuZI3JT6H4eoHH0aN4XNkb5+cRjBJAylw6zXf2hWhqoDbj/pWXlpNiIujakvL
fhMKn87Ma1Q75tUx8XmjUBjTvk7XYrznmE7ZfLQ0gZi9FXw7VYKLRIW5L69tsa5H
ct9YWZaGOduFZgPfoZbQuPoH/EnIOuAo6UqpQBOKURoqwudGbh2VGo0R0zpPU6/s
YRZiNqh3DsYAVhSa6EOodQDzoXp7RmkOwy68RI2DMDeg7+VNM0XJik446gPj6WHD
vs0RmBIv9OqhKgJ6Q+soxp+1U5eOP3PhtNscgFA0Z4wZY00s7rSJ2Mq+QJCNR+/c
1xLGQix4kz/WVWP8FlgtnVKwWUl7PHlWI59yoBZpFmaKRJUJr2164wgWZ3ytCWlw
FtyNto2ncYlp9xiBYtOUAvajGl8Jageyl+VULJvTiM5AAn2vSVKrr4VH3oqDySZx
t5HfU2IHXmop8aBBjGZ3axSvGvgPqDZZ+Ca70XITF4dwmgC4JsLEf7DkODQHDWQI
8VHNFLdzVJskQn9iq2n8+QTLi541LIQFMECT7fMT4Er1nsVhJJRxDW0c9jX5Vik7
dCs6MeSNJcbH7nEqfShfRjYdgw84WVwaveNr2A08X2s/kWrG6SiyHQlB8h+yrBvn
wB4o47d0JH9BYjgqSc89K2bSMU9Uwk1l+fJROkY4KIW3moQJFq3jivkn6pgGD8hV
GLg2QOAR/XUwTWhIFLdizrZG9lPUAQsNqpICBm2OHOpDERb+FrZcVcWog6anu/aZ
NhjwL43xOlM/iet17gvHwVn3cvt2slO7iZfTos0YAcdNyNxISgI1LumclKHSeHIJ
7MvKnac8+bPzWlcpZJqsQXTUpXMrYMkN0iRaU6YnfAbWtgfGtby6aVoxVTu05k4p
lU1jIacnWFUt3CKuhFwtkZyEl1JSSlvCunC/x0tF+goa5oMljsKEwJ4DmlO4Kkkm
9n5IudYJmQ37cegmOE64okiuyBau4EUoQE1/UoG4NlYQHMwW7cTTi50nbv41U5aN
IPu6U520Ig6z5X5l/f3jkUG6ayyIkGbZ3eRIUsEXaXWD5K6EIQ5hdTmfbjWbe8de
YAWB/JD9bFK+LyzVjNg5HfjbjNDyfEBEfOZIWvFLav6g/82vTxBT+GbZYM8MVhcb
YOu8fK5NXnguzJwOsEyqV5VzSeyJCBtwB723KwpMH/kI3JDXuEsKlpW1xLCEySTT
ZO4dqIaoyySxGRWaX2T2Tq4ZiYUb01pGTmNznfvl+T4F9FqNAmOmAInNCBlCpB6b
RkXDX7afCKTQrLpajVP3MOBypidfqoM/0wpH23lh+dYs3204qieplUKj7pmw1BiQ
reILqJQO3G8gLtW1q6Ep9xGQZehFAa1nRgiqYM58yiylb3d2K0bSRkBk6U1niQaP
KsE8UcA4eLdWEYbEdy3ThOeRDCUj7x0xzDIFVM0EmjjfWi1eHiFuhfKo0QirpYQ+
L89ApmawAWI5XTPysSaK8hKUc4ynKL8BcN5stLtcxLImPb3V/C7lN48J1wGb798V
+0rUI2e14cgUlm3CRXM2XPIB61NDFV/HoDxFKYYZr3vAA1U1L4wUxvbMrZ4KspwC
euDtCLIxDSY4B2qStyrXnApN5k6XkZsyYQN7tnl/2WBlKv+gOFA5xsFz1mX0RSiF
XCxGHDQ4pKuYP+Wa6E9WOsKZw+Boscb67kbucQ2gup779yubNa+6Jg2Oc3qFBTtn
Z1zHSN4GDoAo3w/sUCDGipRIahIri+TWRztPgniWBOgJ0LZmT0YNqtrMaQgJgJ7T
hR5t92slr8kTDtDPlMjhby/uX6UQhJqhCsrccONS88TXT7K92saSHBzfvc+nIoZC
gKQ+kI8BDfhUjRWY6lK/m0sjh2hSRvz++oQJ9BOXiftaLdgNczAZ3ETR9wAsIYK/
kFu4tpuuSvKLfaphQWBV6+sq5/dqLpkFO/Pzjji2/9CR0jIhw1Lxx5i8jVBt8Zi9
j0DsXuL/ocLCGFR7NYG4JK/CvX/dIX6O/TTmb4XGqyaWRwoB4TtlWBkLLY+oVVCl
C+98rmHTklinGlP1I/u3f/6TCPUq0y007pPvy76QgdqhJROvqHQ3nJwE/QF2dH07
Haq4EmAZrNvkf8gJogvipbwgleJx6wkgo65rcNKfUlkEBBoLxXX3ek2Epqtgrubq
UgkqrWdFwE3uSMzGHPB6F3zJEU4RSAFke7lKQKpnP36Ru9dS3zBJnILWnnT1tWUM
bmisain1egNwMJkaHm9ZJ2dTNmK4P/DuByyOyA3zau4WiW17bL+EoN5kXUu9OnTl
8hW+tTt3DUbbiPybA1cfDk4ixkHrLlCQOgfYVwHsAY3iraj47r+IiAOeVFbJif3z
ZyOzervWj/Cwi95r+UCs3qk8BTTh1t5qHk0XqgRIeAaCQqkxWWqpPgjayG7lHESc
GJLTMWUM+JVjpGI9B8ln4tjs0oKHgfIztm7aOSgEqE7alm64eIXfqsWrsbaRHFqH
xcnhC4XUqtTfvJosPsgHEFcHaO/l/PzB+OvDyKtx2apN8pAzvJFppcjNPnhc6CQK
36xBaKWxy27huLQTslMEkbig6rUtNVCpkY6yvSC/q7Dqeq8naa0ABQcxlbcO0H2+
NJMLisxmIHKSzJcwSsHx9NJyIKC/4n5/69QtrSVPE8BOZ9Wtqmv8vt6s2dSvwib2
jSXWJn5QZ6RhXCVpGKcjBEImXyHGQaITJIeZ5SYoWdHxj7vUaAXI5wbp+WG4qBcJ
bQRfrTCq6qYyROXZyyhJYTNmXSo+16w6BJFvjpMGizBHO+BSaI6dhKHcfplg/r9/
WtBqgjqCH5OIRVX/Z9fXVrRwhKoT68BlLlu9rW9wCDhGZD3FE9YhYL2R1Y2lYIer
lC9+2ZpbbWqGbZC1tiv9xVr0SjB/Uqd9VdP2QAbFF0ZPKtc9RQWmb1mkEaX4zvS1
rCMTV2cSzby97AQpRZ2ZBnKVK4jE4dh7i8w6VbPMl7K6o3/MIkOye2gJXOCdhtHD
tfI5ljY7arpSOjl2IclvlraZ/4v8uQUNHqvTbs3myTtVtkzPrROUg72f+vCRibIz
ebb2Ukkp9MDhUFPMhUFVOyVZx/IZyyi6Jf7wLI1NXLrygmm7OsAiUkLjDJYAAXkf
COQvBy5WBwil5cJ6VkPL7pgFUzdtRe2uzKPlfaTTLeaMZGhLymF+otP4hB2IzK4n
BLZHdLV2UhzzxHeB4H51HLCA8KU4Ty8b6fyxi1z5cS3PDbF0Hu4GzzLNRedyy54p
+8tSnkgIxO2+3kUptgeNazuSsFLX7wIMoJDlyMt7Xmr3ZQOUz39tlW2wdKBrcuZZ
14vjb/MK5Tde6DmxH3Bw9zjQRyCq1GWp/RE44mP0dZbu3qSpoMM1CIZ45M+i6Tub
KEgltHr8tuZ7sfDLylhiERCvOg+waETR538ZPIU+gfTJHQUlKxw3+uzJ1tNb2VKg
UDNYtLnO01ijhyrj09ocZuJCbHeuDEqaYvvm3sjH7FoSFiEOS9vIJTTeIaLep4F5
8k6YZNKRILykS9ps+DDSzR8K7i5doqCNBVE3fidiTF4LW4ZvwIO3qyNjbOs9BZ7G
I00M7ML0V5qsmMFU8MlNBe1VvJTz1qvExGlbwiN9hPeCxed/kz8cO9N7jS/YtoMu
EpvQsdyVc9lVDdU3Q9zeeDsfY4O7aeqYSgMRYQer+Tx4btqUYc6SX/l52c6MN6z7
Ba4egmBOvE4IEe+F67/fKCL58cxc8xmeC/wAd62M1AFhJLW3g8ML718jEgdfEd88
OkTuEbEz/qtwttebLh14dAZqRdnMEVpsChuFKBKupHod/xRQoF/BmHjH6dVWiJXS
8sjea4rdBRUOrfsuqF8dDgdfvf67zRDnyC3DdZx88TmxTxUQQHuteoQefttnTGa4
gV55uE5z6dc9R+Ur8NaRJWJmUrF4cXfLKNa3otyrb+n8N7RVuD0r87O0L0dHqg4V
sfSs6L2MhJpW/PoQKaYXeRkL8gkAot84NUzH15S+rLEU0vj1K0eeIimaiTyez3tB
hU/ljHN3sB87U2v/QWU0fTTTH+HfWJQgIrScold9OS+LmSvM4MbzD0o05rvwFB2V
MT4PrbLsOB0I8GI23A8SnKysEFVXxAGlXlPqS1mr+9OWN6AUzROCbYW4wXds5tge
R23eD04lVoffsnSBMbhlwxsjiRP4GKK+ZPoIniUvKZNQ/SpeEZrDcgw/78FXSYEI
UbKHsDtWr1D+yxjtMFCZCu0jkFmoHgb4S7laEhDkPG/NR/opsreSZGP5Z5OiGTUr
N4E49oFLUiIeC5hL4ENNJMl8Os4+Ngr6EypsIYsQmVnysl86oZt3M5ZIWrBl1xUQ
i9KX8vsR4yDPJLSmt0Z3ldbaQi2wn7ZolYU5qxd+PyFt/EG9hN6BGkNDTTa6s8Fr
xYlLInDyvAHh5t4rcffQ3FacgREshXV/k0mTM4785g0mfp2vjECMCsnMQy7QnJiV
LnFGQOp6/V5mW58xWeC86+SkbP0R/gagk5A3JZZ61v45S2ARCCEK/cN+5veH06A6
ffnIrUW8a93NnyeDim0GdBTXvcYJN1hCvgNGhRnxiRSJsa0T06YmSl5ggVCNjMZx
lB8qicmD31I76eIqpTbhnDSFmzPiQCt2RN3nSYAMH9Ithb/bI/e+mUEz3O0rEJTG
fVabBR0mC5iDX5Z3L+U7gPOjgKfuc78qghnFooVKpKQygnZoB3yIFEpaXPkXr30f
LUC1X7pWgdUD2aSnavY91ERV6a9U53GttyJQEufEu/8cSWOg7Cp/43QzLnwohH0D
/XoU/4XN2NJSaHQtz7VkPcv92QDO4Ozs+q2r4QgsPeC1UknHgsHvnFNA5et5Q7/O
Ni08iB2j/hyn0Ddhz+SJNS0BD8WQV6j64kdzbvaTQ9cRV6O73OqhiZY89XdPKOhr
TSdie5Q8Fyf+l2oK+BR7b2NIvNic/t7lDdZlFeEf8PQGf5DlbDntjWDQJbrEoJB/
i+2I2YVuDZZPPk2S5GEVYb2IwtYpHMU1HfnmGQbbukGBkPfLFJ0OKU7ZMBJmVqQk
oEN+HhhhzD6qrt2R+i2GsURP2Mpoi7OZZmzxLwgghp9u0t60ESntXzHBY3UYBlAV
F5W2oHwb6kekRS5A6JiNROCBX95t+uvbBo6SyGyXK8oN6k3i6keHrueSQcITe9+6
vHg4aeHtP9QDGtIOyZQs8JTvOw/ipfhKLCT/CJSZVPt2lxdM9wm5M+JFAN2pefAs
S41TVHsvLEu/Su8vZF2y7iwbM3yLn3Zbj4ONu2bI6gzAA0UhkaUldSEoAS45/Pfk
8vPg6PcO+IM627wbewCsADshSHlVSIFHot4sSHz0GBN5fV3GCcqcE6qBnrqS63af
UGINCgvVmAsMEqCaoPd7LVg0QOzthswkbFBPMvcqEDN2WtkjHTufQQayFEyYGpfE
BwkaRDIlLsmu0jYdTFtx2FrVMxLPxkc/sFXDJ++rr+zW8PI/Jei4tgwFr9Kua9Fh
tbWyGEiMlcx5DYzdp71Ku8366H55ayKKwPIlqxjNUTxslHH7QC7Gakszp/1c9Joi
Dlc9f3AaGA+zNyR5WnsQXl/+KAwzoVWfIIf70G31o8iiRjmtac+IxeA4t78oV6Ig
ekVUD2TW68x3uVhcHiQZO4Q7qAHjKS1stIBr7gxYrgjdnrPlapAXsdYpIFDELiPL
ptjoj1S1OYXccQtLIevTExqAgQzsB1nFaH+Wik6ZAXvLAjEVdZwyanQPbufiGUaS
K2Wwyru+bFJhjSoO1IQ4+G4iUuuVA306vDxMjiP3vbLzmKAvhZvn3FIH632BRcB4
xRiWqNeHaA7SPk9E6G8i6OhpOPX9xu7uVziXizb2IaxQQR3kd4excKZXpPusoxBc
SkZHLqCORIf+AOkOt2rGKlE87zAPWMK5KV8YMsWUH+bUU9ILGyPrOpUmI4sltHew
lEXzKLKES50Fc9eEspEmq0eolhbkZKrKdGtVFjw7L7mAybh9HoiwDIeJC1bj27Ao
1UigyAp70koczNLAm7peJwvbP4RItBskCKgenKl4vQKpMtYgCSYLA28qscLpCGyH
sTolQ2qNlmVtu63AjiwD684q/M/h4HXw4pJi+mrRICi4SKeN9QDrFfBYeSEVlndL
S2FhmaJxI7P8GQdMDhZjPK/RFIcI5pDMQvHiTIq8zaffJO/b3+4n6oIBQU8GKmnk
qNZgGPpuKqejOOYg3QpRBOPJ7Am2iV8QM1ptGhWaumNpFnz6c+uilt6HCOMpGAIm
Fwc+niZvNamizttE4pAOhKgSC7doi+VISY+/Uzi/IWfL5AZC1us6Kn8tAeIyc88g
HTF0anf68h54+kxyMUnrQD4nTrxW0xw7nEVB2GulH6TOdYGmBGLQlqjGnKl22Iv7
1Lkb8U7sVRJdbi792tchru1Vu6aPQni9+Dv2j9vi8mNb49FemunCfWcgXu0PWxDx
fZyQHp4GKd+8sWBB3Dn7ecqqc65MdjVx1EM7Vyc0Rhu0thQbl+zFcwYak6RV2nlr
Hila+9HZVEFOOBdC1nyCRUJM8olfXtb2REN6YhtOIiQIr75K/xCQ3gCZYStcBIVp
p1DWVLDdC0EuPT+D5GEkTrCxeqq9Rf0KG4h5KqbM7pm9KlNepQqoO/gE2rZlF5C1
Y6I6jvdQJn+tKEAVHv38BkcZx3kfIBJdYJuin8VLhfHE+bLDE5wL/OEYIfY6r+YI
VDnzQnV1RYWVtxXVfmqnCLuUdMTO7ltFPwARN50VF07Nf1FNIsM+xPp5YrAHStf6
JDWIwAQ8jixMZPkzVufraeRoGCV8Fp7FosgK/WCKEHf0ISxyuUxJ7XF7Dg40Tr/z
uiENPv8URtsE/50lk3qmRq5iPN5IvwlGPuVB8iTi4M9IEHQzqAiTSWnpMGetY1LC
GlO1TyuAXs9Gr3xWFOT7w/D2CK8JBh+BmMm3CZ1SSomtSgIpQZjSq3NZqKRUWttE
ZQvBCA8oTvTPDlKDwUAJ07Z6Qj+6/Uu7PFA2HM8I8ilpSxVtePW7YH1P7oMUcph4
sTs35sHyTKb40SZde4gxbu/I11AkjUp3U4y67A6Tp5nj6OAV/s/TotZwlxkBuHoU
VTSINOQddbmH4kjiwyvuE1AKVd6O/GeR0TXjRol4YIa7YLf441uDpgRVmhaaEd2u
iKD8nGdR9o22TLO6b9c3iBLTo9f0knn1gCSQP9PDw8eex7z3ZIu4Aiacy0z675uD
VHO5Y3oj4xAE2Vy5NsiKshfLfIMFWxzDNH5JUrguQbdiwSMYJhCm5LF3Djd1p0xF
ae7XpBLDmXOU9U6NpIATEuGHXCL1gQXvWwnkia3jAlEL60yGN3wfKrh2VKEpg2xH
BBUrARJEr92MpfYvB9/54F4reQ2Xf5DLgY1ld8upzWT2ZdR6Y0Nb+L4EZLs97qMa
k+pWVYkPKofzo3WdpGR3KMhzoAfGOBRDVowrfh4Lvbw4NhmvGjpGKdUnMIs2Y/Ay
TP5F5dkH3HTb5IHmX3c1jN5hH+T6JNyBH1BMPCclh7hcBRc+ddMQTuWGuS42gBiS
jTHiiBFjIMO5nDjbWc6g9FM2VMQ2A9PTWQbP+fZpCxzTd6eOmCIh/Hr7MX92A1WY
2WoOHHPx6TA1vAR34n+rtbg3nyEEQnRYRBgAjR6AE9qjuCpGd3L1AkPx9NN48sdR
Q6AA7t7pnSaaWNYLWuOQkK9oz09NmU5YKmA+S3wgSrC1MV8RH/k4FDCRKJKOBA/5
wY1L9fNZSAF9k+Z2aSVtNkDwh4oE4wR45YOW5Z+T6l7NYSedcTgRliIskm6f0vD7
vPyVKL4TcypNUMqmKLVK1CrXm9XGY9/YO+WfkbBkuIaTxVi/9OSZLqe+Gutl/BJ2
nw3vYMUeCtO/yMFGL2QfY05zN3S1FuGxR5pCR/xAwbCzKh9fc8N4W3QqIlSpCetH
sKzo1GemaET+l1E3H6dQifQBzmLI1alb5yw0UrPv1gyc3YPHGpcUb0d0w5FYSgEY
+cpU694DNmHsETEpujy92ACg44/Dr65ausU8so5NM90TGOcXvjbEaTmKE16Ax1Wj
HQrVbFBi0t9UCWSem3Tl2BAsZcvMcmsKZ02lfxZRpz6I3vUR4CJ+XzfxwPdyvKmM
ugvY272hkNy59psXjWLg4N7GOkFgrwOeF8UI4dEdiqHxFd2E93iiODnd0oekfGJ+
EY0x2AcYcPrgOOZ3rQXRbQh6HsLnO0PeN2lrfyZlOuWZFCEbdoN84itkeFir6jjw
RRL9Og8RUWcNk5TSwRxM++ZTzBZovMEUqZCXHAxPhpCzgrOf+maBCELhUTNxRl1S
R3kiN0R+W6YCC6osP4LDtQGgM7wC2fc0ZICnyN+tMtpcfEY+SZCKqWlsWtY/dUu0
FnJLcgIiTYzzzK5xCOAZ/7+HEKk+NUOso8WSStrqsBRduixEJOnnvm99ZGzP6/ym
cj6vOTWRv83zXw0YuuNpYYfIfNkdcg5e+a1JXYagHzubE3xTsiqxENaYAwf5dZ7/
K6DoUVtWcbUUGG93nNoMbkD8FQ3yU1wuPUoCS+GRwlnRdm03d5Ekzfl/KtwUWPh7
ihr5WQkxG6IsPMfvbq7xl3Ve+E9KC5Ia+JNC+X9ev0rb02MGL7I59UbARFTzGvLm
NDjTmvz/kSVTXna1LmTQBE7IRYnhmAXDVNShX/y2/MXmNtPGRN5OTP2NbsZMu3CX
8373RiqLPWjj7cvLOb8U2XoM6O7fPYAC/IzKPDDSr7Gits8YS+V2R1qjq4YIb3/p
oInopwfHuw4WMf2+h3V3dblmL81RPnhrYE8RiaRQh3kFegmRp8SuHHo71F17Rrre
OyndTe7FjhtG1Q0rk5iZvMQTZa55eGD8jK2ZNR7cx5m64iVnZeEsrkw101dPz6Tu
8RRD0V4E5boYUPP2eVb1AWwJIgh8yPewhy+p2eKEoComKx9S78afyoj1cWngXlyp
FGtJCcOybpflyT+gctdXSE70M6nNdVINvl/G8Y6sc/6q6+DeCGtM/fIq9sEZa2U9
+VCsOxm+4Il/zq+o60LSwHuUEcF4XAKTXSglW9hYpzMELoc1hC4SKL6Y0pIhrdhG
1JvS0CRz6T7Ib+gwB+cCRnUvxT7uf4+ufZ6fj0oO2hdaEGpxr1J5gQyI1MgB9S3n
g+TpNCVOJdWvCUtbQV9vgcrOwit2OUTLgDs6IqbrZV9CWyUWWOIdEOyojuIdZRFN
R+NnLf//0icrbLzCsjWo4nbSeGXtJ6uL/JXeddhJpCOdQ7U/NctFPawD/bYmtDH/
6X90GOg9uFNWmT/6k2tC++9r5qcEpRDccMIeFWOo44n8jruEmHc3uUGSgfYSJ7U/
hyO7pBGfB7gFX+k5CLu6n+DXdgO/2UmJTisjsffLI+pphVVDYUgk4Ku09/oHP+yh
gSIxTTZ38Xn+ULczyeUfhCr0XkkUQS00AzzHJW/L9Z45YPuD5PpSddUosomOuLhx
8jNNB3248CU1inSJCr9YkkPx2E6Lw6KJGE679cX7SIdjKck6OYxIj7N4s3ik3S+/
XkhXQ8yge4FGcKrDBIzXIqjDDuc94RbwArPWOyJmf9Qv4StM5grAeSO6tq/xwI1i
BmjKMGZuJf0WxUyAy9TCa107hKh/q/LR0ZhtUPo4bfKpVXmDqVCdJhP8mDoOKvK0
/VcDdssI8fA7jSRUrO/AvmPSiqG/Mhxpf5L93e+cPB8GKlg2s9MwtJWGr2Tr8IXx
DM+AFLgpOycHcR+wjLiZm73ZXD10zs+7Ez+c1k/DxxhX+g4PA9Nc2qnSmz6+EoBd
rKjkmUEdUKQMK5XPsRPEM4J/mZe9gVCcqT0JvlgsRS0g7zgDC3IWw1UJcW1JMTY6
hTxpMqMpIuSh1SKP0Gjr+789OAIDFor2NvCswThryvJQTMF7tNhoN3wEu4A04xKe
BT3ENBq+1uLRwqNbt8GqbvgOq/MRhmMMysNaWmmYplcHOBcDrdbXdI37oDSOLsaY
m6c6jefFjZN3hjZh8vjjA5H9vHLxc/jtnfz9/CY9UUMTxgS4tBiwF5Y8WdeCycgF
Dt8t3CDOcUshwXpazPOE+jmYADnZjnDFh+u+tdZezGvkTvd8Z6R2XauoepYJ1M7U
hgdXHLm+LX07vNq/srCa/kOGUc/YvflTDPpZ45fNW43g5yjeODFPfAjyoAa+N322
KEmaUydxu5hc3EaSBx5rVaFnuIHaR8LMglzgXENDwjROxU4zMhyNBm5HcbN8rbDK
YankZwFGw5v5y1sS2yhzRSEA29XgqSjWHVbm9UKcNhGBzJJQFlrRXtQoYWYxtCII
9DgzLe08q7uS5hbUlulDvgTnNQ5dW4PFCmIaCHe0MVMFDC+BguHVGEYYnmBNnTXm
Na4FbmKFxoFtMnLth8sDuW/q+Lutj5SB56d8CBONVnBDnuvE3N7PVsp+QKq71aFx
tybQv7qFFn7YLW3quWM7kqH2BbwC5BaUftX1J9QShZvcyhI5DI0BEa4h1qzn7K4o
CQlAIioH201NFF1iuOc8vBLVBl8KjByBrkuSMxp+7/2g5bzvEPiCTrgVw1fXBm07
nVlRPNvfpfsz/pf8zqnGM4MU1hJRNnzlKEVgCeBG3B27mrcSuL/AgrV3oI4jJRc9
yoz39emfaJ/FLEj7V8K9aT1WHhvh+HaRUS5yd2koIwlZgD9aKnll/fvaVBg8w+q0
IA4XhoWFbAtTTVJRv5F5C4i8wZIeTmBVIA9owQLflk0OO1XQtQEuetytMTLensAz
UsDbL+1C8VFRwkKxl1Cv2FgjtvbJNEWXqUq/IcVk/9pICPZbB6OPxGEYGz/vfW7h
fJaMUIVe8pjs7kkR4Ty09FEyeuP/vREdUosEPVm70v4ygjLuWj62SsGldVmZ5rR7
juC/m/+E+eV336XOJH1epsEQyT0AtdBQHsa7M8bll70udGSh9vjZB4150DuY8ml+
Wl/bear9nKGVLLSJbKcvbxUG0uO78L/PcXhk1AXqQXKoAVP7tlXkDFk/+mxzacgH
jO4YgGit3SBFzTNIr2h5EQ1RQT+/2ZO+rr0PxSPo5JhhBUFnLGz96iImUcj3/C02
clqLTyPQNgbjsB65oenlRrRyMhzI8MGcL+SUjAQUJymLJerkY6JxmKQWeSgeuHlA
RoTy3qsUR/gCiTObETg0+h33lwliHIWhMu9e8t9B9oy2tfvN51nXCZcwqzGVH9UM
FfTEzyyUCjXZgRj4r14JrvRpv7BjUCMEa+iMo0W8d7ae7H2uSA0LThpsyQomec3S
Yx6TWzg3HHsA9TzjwimMvxbZIEKIr9XC+7TjmCSyGOvLwEJ+ErcAqe9ndsj9v6Wo
qjBs53O16ovPeGIANcVDOO7pD8ykh+bxvFEna3hUmE+Db7/hKk1RRmIDxNE5QIcg
xEyuHtO/QTiXuIgYNRV+B61e7PPtvg0/5kksDq3xY9MdsaHIkIDuoE9T5O1uYxjX
1mv/dJeF77aKgepu7cc5Y5o5DKG03CpOBuZMHE9jL/nlyG/IxlolWeM1wxbORpWE
6aqO7WziaUj8xEY4ZwqqkZ/RJ0RxAl4kegux4r/Jr/3xgo2DKOpFj9iLfY5uWthn
NHzYVG6ShfHA7cgGBrMp4o8LRhiq03sG1zgqj1xgkDg2Pv+YG1kyG0rdwxr3AlSF
QSFEpm3B7kUh9AU+ubCK2uPIVVp2+lAa0wSWS9CRQLlXWUEoj8y2VvsQxtJan3cT
WaafZJdf9hdV5FhoDZG9D1T18ATJPqRUGTHWt6AzO/dd9MS3FyOhP76J/ZuC8cqv
CURtel9aVkljiUgFCoownlHT80Gcl4ybbdzRk65JQLUs6EfQyTcGcOrVeMwEd+SS
wmtPqqq5/Sk0tW0DOZQhxhLlrvdv8YEV6ARiiK35FxyXzbGHuLTPco70r0c8epu5
t7EO2aiSY38kw9f2M/JWgMIF3WoVLugefmgYbLz2pSPSQv+GnZ5G7rfzecIwodTe
nnLSt3+Bl0GVXBVgb/ibi4FJGcq6NMsRe0EvOcDpXfrcfKTa8tbIztx7//fptbaK
gkv/IL6sxKyUUzr2RtAw4GT03RSSgb0fcyA7SjulE8RyAOKC+dFaJqoegte3pAWL
ig0uLuqoQWFbNo4z0KFF7nlE5E/72iSHQlH5DM0evIywk18VvWrt7LE38cIRSYxm
dyfq7wzCwg51e867W55Xzuk4yeevonm7fX7ixlqIP59h9dHJpQwjt5nimjY1nXcI
JnUwebSw6HORRU4bFSAowlDXUHo68i55tfLPaIyguUc9bgsZ+dWD2ztolClavLlw
oBBZIjgCjekwBqfJ+itvNGWcmJr5QfXWT+Ce53zia7Sh7oDgow1ryQdJxePUExJO
ZBQLZP6Qfua5b+//TvoE5sWkXBY7MqrKcc5qfSecmwBk5ULYOllhjHJ+4tM9AF+P
h4ohK6wZSV2/aSgHYny29QegbWfCok/d/fXSOuRFXDjRpwFeElt8hjAVW8DKLdni
4PLzklXues3x2AvtEJKCFURTU3UFzLbwrSXBKZg+kcAtmJ+Vp0VKWdJIrykFkCmr
vE4Il+i2BtOchdf5AeEiSHxxYNWJh57Q9ouw6dpavDGGb2xVMGcZnSrzlOw0Ihb3
BPL4Tg2J8oB6AX9bOFdJupYqeAkuNmQGuSxtnpUokGk/t+e6x/5EN/Q5vGrtTgEc
ISvToWv8YhRo5AlrTX75uotLSPI/Fv8yE8D76jALNlUvjjUVrw95YB5T/B71WyOR
zWNnTJoQUfi0ojqoOV8FxdjewNfdiyTzDL83rzqS2vuVoAMQoRwQLytM83pEBxep
HUvQQfCsQpBAXOJkwXx9vAeDzpQTp5C+Z81jXTsTfugGRfNHqLcISKuPCd9ocCJp
fBoGiCVCa0zyAzPB9R8BmikweA+HCD8Hh3l9T0KqRFBPtN9dW3z3X2rt8jgeOm6w
RH6gTmfxEG8yCY4YnKQloZLnt4pQinxAo3PVav0dR+c7ksnkTOPmDcJZK8hzJVEq
CW3d7eyWHzhbeGtsV8waWosyCM6ofHmBddcoFGthQiv3T4I0+YKso8+CKf8SpmJT
yn0wGEWaakc8l0pjj0ewTj8R9h20BD8X3MxFRAOfkeC6Sn1P6KJD85DAEtNUd1tb
At1z807tE4JL/U0iTMWv1e/WWoo240CtLC/4iDqsz0bw9089HudsWs+ACe+3I/dQ
kRZChSACJYrc0im9ef0HR/jqN4w4C/oWAXCyTWA6ocFKqRlYR6gsB6dSj0OT8Tnx
rSIbhWMZozdwYWrkTvMz9Pk6k0f8o922JCTop+FRXWxyY7tC71wK3XB+OoYYdo9C
LeA3T5XCDsqWIP8DlxpmDlkD2S0S83yEQx4iIgFVI+E1GuYemd5q9HV4K/zsD8In
8rO/gLflxjOQpybFqGbngSq9cfmBq/PdjwImqjD9eTwfpUjCFF3VfE5XpNuPQNsf
Kp9t1H02WzNz9Td5uJl7sWEtx7H99ca5uM0SnfZjj8+5qAo5mDwyPy9IDml024hV
uoLUAqIUvIMLpIHybhEaZETCua+pAcKKaEJoWJS/jT+2J/5hFOOLs8W1MaZbUe9I
Rid12V/d3xFu3oUFpwMMZZzhIemtvv/FHMyebJSuXd8x+O+xP4Dd5eDY5bIUfbHh
i39b4SNmHIFmzA8THYgkmWuOhNjuoiWpwlwq84xvih94ww9k76H5L+IbdkcZ3k+D
w7JznM8lqlwZH9XOsIAobCuBTkangq3D8OHMjTGexPIDgJTBp7qdzWVhLZo8c6f6
RKe4BUnpHpNzOsFa0GarY1ybnMJz5LyIHAz8BckdW/p1DuFfoEhBlroBYtSeG5ib
r3W7XPzWPhntBfPL0yFKrFlJzvLeqoSjmeP3xdLdMlAil5KqEiTbU3qapY6bxbs1
26d8nqwoc5UVElHOVWBEwo4rNTQDdGMWdmjjuYTJ2ZB+u++31pJjMBdQNmnXr8NX
toxs799Yacg2yLWJGiQrE73vr4AecTYYhh7Vq7kzEwoyN55ncWXcw57N/5XNgFPg
Mw8e9zEq68XkMtgEnInwUF3GXr9G98xNK8N4i3Fju5JCFEJBU2Xg3hK62PmNe0KV
BkBsIkpvKhWwWt6XgVsV6NHnQU6STzq2vtm7154MX6azW/up9lAu8YVU/Shfl4aC
bnIERAfFWnjA2SwDlU0DAjKo30notypVuQFc22VPsAbtMSnERRD0BtUtULYkRXi2
nF9wGAz2NsnBN6Wzr3ZlGgOIWTH4OwEYNztO0RVih27CNDsbcpFEFLlQzjPEL7R8
kc0yAX1sKnZ+jkIk3iCIUmCN6zmJ96fKRlzj3dmJA9y/76DKEqRJimOx2jEVrLTe
ZQPZZpo2GB/y1TLo/4AGlv+s2ytcirv2mzpHTriUKfNxVgGe8k0W2bOCV5A6hz2H
/t9TQVb5AdzosLfrM105gcHT6tUppPVMVGoKh3K8h3vH/Nb2T1zKbgrdCs8YzHZS
lnAlqN/MR0qkTW0xZRAqPuJFsJmWruVYjCohK74/vZn9Qsl/DpwB+cAx6H+UqjFF
GhSZ3oBAhR4R5HX8NPvuzdgIqFiuv4x+T2/9EEfZGUYVBfqz1t7hk/VOfR6g5+bk
i5yqIGJ6aY7sEHFHqfjOAbgwRZGO5f/mKLkgbVCKBdquYYnjrpjXYLgxLVuZeGcx
+Z82loPqe1Yu0AV5AKNiSewnYiQrUXkFIybbNvxhgE2wWVfuw2EFDODBZ6kRhStH
1P3eu8j/d7QT63Rt1X8Tg2d611hNJS4o6iWzRLlwcevcCMhZw7o/8akdFAcXhyfT
mvs/nGqzpryRxHjYNzGGI3Yft3YhMl+icE1qQtXje2bITjT9i4q8lDLk5AFdAOQG
et69ww7JicyBHe8vhkJUCGICn2H4tOQyiCv7+RWrGkP4kukQmyyYlNH41666j9t2
nXynS+8+Mw1bUw+l7Sj+wmxAkzs+26vLkzL/OFyFiHIu64BV6nuBG0oG60t2l7jE
qVC6EDW80kzmm9qMfKfVIs94w7Ch/l+Kn6V5Ynu/oEDZchyvutfwGC6FmdxbTl34
EyrxZ8ZKoFqUM0ydPI4lPQYU6ElxyeQjCuLwlgFSbsUu99EUwCCr3oDuNpbouORg
9kZa6NjW6HKeXYgvCdPkr2jDr+Fq8UyQXL/ADpWMseCDO1Xi8gn3dRzTyD925heq
vUA0Np5biuYPiDHd8pwZs+1jVA1/85Z0ja3qMM0BTy6Q2wrhcn8kTDPdhYykSZjS
nAUy/177HW12+xpumw4MqO6qXXXVbX7gk8qKSd7BC/6PjBgTEVYH4nWWhNwtkss6
KATW7Ix3XAst/PDGujq+PEgNDVZpsb9mbKiJbUHUDhoA+JrM66gXEwbcGGmJvxiN
Un0a9sfEYOaR1JY6lRO1viCrffmC8KMuN9tX/RchNozGikOa3RkJwokx1Z+VWaPV
DmF+vpdjRpF4h1pzseFCsUZCZA0vNrgB4KjS1OvkLggsf+W8Owf7ad/LaVhVrru2
wgT4shwcp8OID9CfCCz6g2/c78Iz8uy7uHN+AKobuiNYm6745gOapgczy9wTCbv/
aGSzNIjZn40fgZ20ngoNbTj3+wBjNrW8SojFP1H0Lz10RwTkFGMrOsmioein41B7
Yv4Gtm6YNK+KH//VcGo8A1z9hLCDCC+RWL3YrNf7U9HXX0oyisnRZZvVZeppvwEc
X1NedceaNiM/rBxC4nL2ZchBvgcnigRBKs76FsNtd9l7fYFrfDtwd79VjGW2f24h
4hYl+y1j8O1dTsGQIu7h/Re6SoEs95bU6EbqgjEJZjSeDyhOiHUs9FYZhSJ4BSvc
+Dfs/wPUcYA2hL8Zj46ccx8yXx2sqMcpCC0sIQb16Gz/Aw4FDFTDBW+bFcgERFY/
3DXkV7G29jak69utrc62l5b6L+nJ6gndD+gsHKV1ojjKDb//igdWQ44+s5JvXh/c
owjyRkpW2xTD3WMjRvEHfmEywk8qpnWswrM66vo/0UK0jyEuDq1hmM8o57S1OnSs
G3AygK0w7+KnazLk1azF5oRBlODuWway3zIyODq9snC2506OawEtwkAQ74L9FBF/
tSiRzarwXT9JgRCsDsbmMAaWjuV6wNgvVHbVtooHg7EimIpmFyBQoURRLWxzqihj
9DeI+Vqx+M9OKoTLNtbiCKjsR2xqF6FK6C6JtuJV1r0ebhrCJHRCOmNNgJBb6Aiy
zQP+du+GYlZpWAdPuS1E7swPMsk8MyoqTS7h0Xwa1nVAITt9EA5REyV8em0vsQTW
FKzp+yXA6tC4h1gloh1fLTnIKuIBeD1LHebjbUBJVDIum09zHP5M9e9ZaNGUgHAl
phKGyFho2TIMk7QJ+o9crS1uyFn/lzJO9WkVKMSZZXe1/iVkQKQuE+XTEOkkMWJo
rBXmfHU1JtZLaBDSDs3wO0NwnP5nPQHdBmtSVcDeU42raGJjLNfvNHOnxRFgDgx6
Qaa03Yzp393+0TRLox/hj5bOjTFWFiCPLdhBPEokGdB8Dn6xh+J7C2XiwClW/+Kl
Ck1v05mjeQeqkrmOU5aVBgx8vXocIDNab+SxU5ji9iFKGHWPSMBTY2lVkOvDcfl2
cyujwdlmgH9vGN7VLg/nw+my0s7KghXn0L5YHwQJY2uNdd1JLj5DulhL5ELiFpOt
IUWRpMDCbw1zpzfwoo6j3ZxGHZOIbETDbLDWs3XsSrAl/6HvUhQZO8m0KHPi6q5z
HPsH5BOxDBAUFOaVuVLc9Pwd1upTtHAnrSElVesO2SfujeSiJ1OPu2OiHq+DZZDJ
Yle45byUQcyTOiSMYD/GOlTBd0qZY2TnKAIqu64Z9wmXlHcdtAPNVob23nEXaDYu
VRLeuE8jDHlX/ukRQusWNWvNfJddDEDFcaElJAeJN4xWhyaUzZBZBf3LbkCUD7cH
pfGL+p3msXHq7ZFi00JuVrzqKHAJRjsPfWmy5+40JHZPFQYNajoyXWpWOPeAtQEz
vMOFSagl7L6PqX/yFFvZCAwl2YO2FTeUcSGl89JQlMnnXgv0uUk3aw2ZJ8ih/kSq
//4b1nbkHtB0OQ8junUoWC+TosuPa/taIEPMaTjT/kZ+JTTruxdVI59sQPKhrysU
HD9KzY6G9l1PkQlV57oBuNnHPEASMjnh7g3gKHOiylNDjKxMxVr3kMl5teS2G6TW
YEuo3+ZjDPsgMrcNAG7ZEHtX2UrVk+RIOJnC5iKrR22IYXinGpdYdwuv42hikQr5
bEgXaLlGOgYLCddKHzYCFsFck9LraJOZkpVYzDedzvhu2zuL+IgfyKRBYu6R8Tsz
Az+P9k7+BphgVjqvBcAuq6seSqrzgwiCtVUfhjgkd4df/7VwYGDrHC398YFr72MA
1q9C4i2+4bf1exGZYL8IM/yl3VmKLDcTTtiexgXa3iRsJwvwfQobbLNL7elgxNta
/f52f7yTfd8VSPC6UuM4AgU24LRWAJnpznpGemi+Ge+KcWpClEYAKlzuNzRVoN7f
/BylVGyDboMVHMz796ipS+C1dr1x7Lr6ZwkqtVqVvL1RYTjcg5eg1jxzXXb30zKv
SS3r6fyArG3iV8kRx+XXroa1oCQ/c8mmRdMc5DBrkLRFC1txOGgs6nfzduIa+B4R
g+zNlk+wDZ07NvVRap4mCQX7OgcVglkfcmUtb1h3xF8LYkerjU9upXBc6qjUzkmR
NeBNAoFftm63zCgeQm6399aWERhD/bS0Eqluri6LlvIsct2KSGvnH4GB/MfGxLw+
kSZPYczuVpzqAE1e5d9eoCZPKvKXd3SR7cAUdiYXVeokTa+tY33WJgHpTp56gf7F
6HbP5402FguYTzN5lFSXPeB7Rq3E0aQQL6lHHLrPOCpc3EAR8+lV12wW4HsGZR6D
8xjObXRPIs2ZlpHQx0T64VcrzHFxUerC11xLPQNnhzoHZrM5kih6+q5ni5oXIeIy
PeGVKcPxtIadaHrqV9tl14PSrGI/BsXWrhNYH+0eI21pdLkww6+54FvN3t0IYqG+
BHsbKpFyFjT3eIuMhp4Ilmg06Qavg11zy12arGZOpsq4YQ+WS4eBPwm5hIFsxjDn
gJ6271evhAVAUwAiR1kxyjaZQv3FqmqCZjK414OT4h5bHsmmwqrmUQ+5Gmam1WDT
KRnzVPPmF1QI+bozhZsF9a83if3HIYyslF0D3mTI7PPZT+RbSxPl/chfkqa4flHS
BdeDNPJzTyR6eAWKOwleLwbZqk9LaB+uCJ/AgUGhWE/yexf/feUiu0OAMNYtPyi1
aghy7vePqGU4l3lsj4y17JtwEM9gcBacGr7yIC8bhjUJuQYjv86UVR4xk5eGHjLU
2vmhhZmX6cVnQeFNhBZK+a1lWs3rCeZEZ/39f4BHoaAucUnFdHhRO35frFFSrI9c
eFXuSfsE6zYAjatkqcf4DBEy+5csqezkfy+X7JP4t5EvZ8bMVuy8nZFDcKKBPStd
BhDs7LgS2n2V1DQ4dIQ1JPvMTa8P2L+eMRUltxQ1iJl2eRcc5UXZzs1vWML3taqm
1vEpMvxTeXpyNfhvJNAk9B5QzU07JVNdS9bCVd4BvqQR2Ma/ISgcnxP8Y8Ilq5EV
E+LMyf1GEXItN/QYZmmmXT2Vqb+S8sCgjZCPqfvlVdDsGzdH0jPVhhNCKwzL/eij
6le8nW67jEzhnLxm23T9kgsXdr792qVbfemddrbdeqgclo7YsQP31A5uzmdouSnk
Np50DXUFNee4WYgBvwQN96IJwZAdp0tgJrBOlsCe1Uy6GpGjBGYKZ1Lc/4SDG2X+
uUOEKoAK2xQ5i1u/z4MyJJjO/9opcXtC0pP4GMkB7oVwAl3A/5ohN372fVulqOAx
iXY4x3ysDP8kQXvqOYQL9NjE2Xq6XyPGYfdCTmDRw/Mww+n5RsApMukNECMwOrke
eBpbpx4e/KOHC4OqgohLDuQkvDyYQGPs87mX0kTycWOXF5Cj144Z8yPzTKKTLRqg
JMz/4cuR17Ou4hw+yDbwS9A1CdJEayvlfiF4/MMrT1sWu9sjvaZHAw6k4/jZGA8Q
I07KmQJiG8iroRQDcVWw1l+9+V5b+8WOVixlt0X4fOt3jj/JcvDBnINCaPQbe/4Z
dxKVW2o3cxMv8BWd+fKubtfjfpjYcpoGDsFYKgtCI2ctwUW3UpxYxG/YBWvOY+xZ
d0RmepKWhCy/EVUz+qPVNNGs+8t4DLAwF9xAPZEnottU9S7xCA2ortQkj6mXvwYB
xoADCmgUKGrXQh/2bgS8bzEGjnPpFHTc7wl4u0e1tN5JfAyZ19JSzBz7BcFE2qpQ
jqfb3nxxgdPH57s5yIwFwScFOFLzLNcB0jsYnkxso0DBoxPYeQg+FzmEmZ6bmEwv
XnVjPb0nvRWPbOnC3eATNYue/BsOHZKLTzWvB1pinIfRfNCEmfehmWSsnz7LrVQn
WVYeS/Pqz7IyZ1SlfMzPlG9m0XNqwUoDf6wU6vZ2H2wDulBOGHvuOS+OizqIfzg+
f/pVn295w7OGLzdrvH6uPu9HZLZ70UNZ7lGnYgvaSUAplyODhoYBrRWjy7R1Jk4y
k/dyGQrrFqtUFoGnJdVH3bJY76Q62tbYs9qUQsIK4R8u/EOc+8kIkPEKBXctqIS2
fUA7DqDds/VS2oh/6E30WoA9dE8pMPuLySSGijwmtNTOqr6lqafhs7NcPb8786PF
DeT83CNR8l+V5dTCqBeKkJYotRpihSQe50+59bti+tNWpzZPi4TndA7No5DqaZ1d
0inOJPte1fZlQrfadzoutyDL59iO25kQHbC4Q+CCHsQ5iqVPS4CTCpC5eS9NKXZg
YAE23C1rJtKgF1o4d9JJqT/cdJz59yfiFeLc0ednqnZ9uDEFELG5LqlAc9H1TkoA
SdvrVoeejxEYUh6Nfwsl56H1NXlOms3NURJPz0kz2GvL8TGVV/1CVTLP51Ra8ivp
NMHa2qd6ZYHEMSSvVIIqvxQekgVKHgzTf/gaom2UbymT/dP7cUuyusUnbt/ZfUQ8
/t1caDkOBEqqtILUo0rUMtuyhbYlmSyVjIeqpQCCL+87nd91kiIQT11Uyhbp6nYH
xqxtJvloVAoeT0RJ3e9IZAvl2lbxvjUHP6SHt55kdPkN/gp8JDbTNiOgTSh0q3ne
lIWXdfptzPJdZngxeQMwjjMXB5ybY8XHwOwRk+06cuF2tikYprZ0KmyUZ97kFyz+
XsvY5oxMVN+3rPsSyu+XzsBDcLBQqyWiR3lSzjiLiNtj9sI5q76CZid367KLVuQu
8hPvZwqNp4+DnVsHCWf/D2jYWf6qT1fw/fi3RNYJrQGQS6CoBGz4zmRnqW+KdHGV
0r29xdXnS1ud/USokzcTGfT6bml4Y9TpY66rI8h+rZ5uc1dvQnSZS6fwOLFH907l
Qy/dD6cbPNt3IBC5EM2CX9sVGIoSAk6zVBwoTXvY3fReoq0B0i6TTrG6LrRYcy0i
lyvdTRRhF+mGqhplhYtw1l/5jyl4K0z45sbmwLZBoaKAiNwL+EqZGvRCGcNr/Ug1
8zG4ZpXcpu0YzUIwtiUyHb4B6ZGe7LtPJDDeUlZvsJsz9wp1XemG18XfYqwtOsdB
K5N0GihMxXCZ/UGbMpdQUAeC7WTeZAUoG6dC0HY3SEh7tVrfAgh9ERtM5jm3L0Ay
Xh7Mj+jUgplyQH+g/CpTWMBuX84hFH6M30e47AoT7JNBpsmQGM9z/Q8ZSTQk7Qdn
Eh7z+vyWkg0iwnx7Z/nEPVpClecGIqV1op3DGO2s60/M2OP1+cY6btEV51DzGq6Y
3y3W07sKjVWWU7jUNqWXEqxwVgmIEGFOxs+yw0T7nQPhPaScF7VrGn80UVIkZVyZ
CPUvjUxCkjyH+YX8VZzpA0E/H/U70nS7z6P94m+oCEzxkvkBtvdNqnZPFWIudb31
L+14Zh7pldctPlc6SZMrtlM/UE0EL+6iQthnTtBTSB93lOQmpzOd7OECmiG2ggfP
p0OUzhuOtVLoWJTkl/lVTJvSNKcDGE7ReBl1DlhcSGwwbtsTiA+D7d83TJmPOkUT
KGcGknSONoozxFPB5+NXy5ulknL8bIh3BLCA9Dub7bLnCDcm8W1+D20w00uePk0u
+j2SXLCwxvup3ESijgassQb5r07k9QDbGZZ4q0HvG0j7+WJrXw4lfoxHamKty9jR
c6hXfYtXScz3mxPA2fPbGRmK1c6UoJHsDTtiluJHpo7sUtAXmH/QSCioTn8x6ZoB
JIQcnxjF1pUpxvo8jyX6ALB7269EKFtmELO/PMUSrEnJduDD7Gjzri561sY0FBKf
btW6u16nFjgMez+b48G16JvIzkUYXbG9fUuZcbU+Yi2q9p39FoJG9NKb6inBpvHB
YDjikyBnKBXyhB83bjNO/FO4OpGdNdU0+mmMyoeEDsmLxohTTbXEMFz6LwGxLPr5
43E1FiR7d8msocbiBrQIzztxNK94rypvrRtZfIXpdWLyI0X2Xzl0aDl8Q4ND1nXq
+L8MaqeleWsQQ4I/YdC+vnPp71+O5PUn614rfmwPvJzvAmqzn7BcRoWzXZN6rA+K
k4z7NxJ5hnhpRqObnBI4kp+MuzITLYw6qpc+BnxbmOQwSjNxap0w+kkKA5zIyufv
Rn8+pUHlERWiSAcE8lAzdc0qeL98hfhjpamTbOUFAddnv3Zx8I75nRaAza9OycLq
teG7JLCKUEKBd2j8j1828pNR0HRS7LT0mrAMpMXxSal4IZqSHc5sJMnNQ+H0rVDZ
gXc1CkcW+cv3DNS6nIHMvQ3UF4NbPUO24tpJQ2l4HPLFvtFea8gaHj9NVa6hqklW
dqLC9fDwuMt3DDgvufRCBE7W8w+urv6aBUt5HQcasj/MIEhfw7L6qUI2uxGWH+X7
CdP72fTpO0PyCFhibtKldUuq0f9kxHXZKEwIYWPXwyStLaJ1zwG9QrXPYRsVorMA
zoQ5FJqOdjMupeWOoN5FiD3hWgAhqSENtXM+iWFjkgvn2RHpAQNAwAXgseE+L9ax
Ti4M6Rdhsxu6edq0HmPukfORTIBW7JQLMxIBgcTfZ1T/Ehxd3Apd7Mfg2BUTI5CO
O6+L5IlnJU51iIPWdSizMcD/+COf5GZFKgqpebusRIBFfFzH6Ok4QnJXtwBIZZ44
Yw3lUHXL7buP9Sgz44AZRKsvPkaFwCN5Vund9j37RMdPQyaHrrImLvFOFhjov1RU
N9LQstHW9mNcDEBhyMLzrN1orUuyvG9sYnWbfBo8rOk9kWgxj3bIbVXA8Q8+bJPo
H+1EKeqFzo2hwvQUxx3g001/32uJ9NVhdCEG2qExZoM0T2qk7DGO8sbzuKu/krUj
WDGjnma/ngrbBs6oLP8pl8TxSIOUHqiTTg65db+7TCKRvq85M6Wqq0BLqL1T1WxS
WtDDcLkoqzxPgBxTFPuT59nSo7CjKWqT/b4qMSh4Ws/XDkvkaGpUqyEhw9pqy6hx
kvJRGHL5db5rRWmrZU0bGayIbxNXo+f6a+/qlNjd/67ZBiAWVtK+MjM7tp0zS7fH
Iv0xqKl8kv9iMGu8woaPwtZAc4Tg+MmeWrqa/hvkHlB8+RGIkXLPgqeUI3mXmaaM
/aX0eIjvgMd9LyaGyT2gqqQTKjGYr4K6sC0fMeO0Yru7tt/dNxtDj3NIFYZfv6rJ
jNONFZl89zhYLteU8Hoye8nUEB4pEI6OpSCOiFJZ+Nve/E+8KNXTJwpP0L6cdQfK
rVd+1r+Wl1is4FR8GjM2MaUFMeTt9Qw3grwaNpU/qqpHBjmAxh1GkvUuhYoUmUda
12TxcRfBE3pyRFjeeaH7Xn7tKYWzjV2n0gt5f/iXA0s3U9cOyFNeTnYTlCCs6mTG
whKuIk2yJ/e3s39LqJd2IAJzm7HtvcRrSAEWL4FuROwbih+Agn5UHGIurw/QrElU
JALhA/pCaVrmwc1cVOw0KROwsyI58EDaUZ2zc6WPhjDIMMRQev4OoK4rhbgVWATg
wIKwskRs0RPk8WsfiNG3I4HnQoWcOACzsuv813abDT76ToQjSEONlo91L/yXyNE+
ZUN+AapFE6Xp8ZACVeYMg4+GLid2kyDN6LtCb/QtIK2eXV1o/ovQWbESj50DW9FR
Gzi9uQkVUs7hdrGZ1E5SbdKaygyEmweFwu2tpO1MAnodj8I2pVSG367RyQvef2jU
PjzHoGUAjLiWL1xo8vNMUtToOna2PtTLSyOhn7uvjcr75Ft2V1CElg8irZBEMD/a
OwwTajooBUHJqISGw6Z+LSTuY70VJGdZhTZ3JjfmXDoXeACVHuCYp9dTV+Vz+x75
bus65VLRkoStUGOBEfFGQeb6JTI4HSfRUu9UvLDrb9B36eHZsRTO/zilUgPSv7wV
PWDlaaRQ1z6zhnMOeDyWzAlObDwYYEruvaq66Cr5m0kIldL1SCT/LkZ3hJK6nEiU
GkLugJbh33gr5DXyP/7xDscKJsQkIz6zkr960FUbvrijNCIR/ZVDaReJBn58AbNE
36E6yAV1cHPDmzd9bhwGGLlwyjsc20Dzaj8RZzulA+SFnpWiTdRq5yFzX1n2wic3
hRF2jtI8WRnF1GjRnaCJiX57Q9NsAB+mUfwzlvnsBm1irMeLd0kkjaVXiNoArj0O
KTBhIxFfPmMR54d0x2k01UA/mi3xEy8MMVpMJ00u5+JWpc3Cq+jLWkKlDQ7swrCO
gPgqU6FNVYXR9uujb3rCCowcBnSV7HwV8DZ90wFSf99UxhR2OmBmdRyjlavtXiG2
PuN8thZ/pnkIK2aan0DZ0MrpdbdkhRcQIfhEAim2bq8+Glm9FI+Yo9BiytWAjHgD
Pq9LjCWlw0W6NpJLGAVOxIoXDwUx6Tlr+NgIaBJmcDfuUX2xWYfvHdL5EaCacyFH
XElmcx3dPriLkTJ8t27MIoZ/xJCOC0Dit3A8V6yxHukIn/jhMY5AvY4EJol3ukKk
kUyen1z3n0LF705Icl9yZcNJIxcdSa9BcnUzpkA2LrX7Dw/gGbB841PRbhe0mbeX
Fu9ruo477nDCQsE+EzIjoiJwqmJs7m0fukHFLqcZdh4fOI0J922pPYmHOVIXdrLC
sUvgizmL8g1hkEYdFlDZbykbm8SQAzq+0/VklYM/qahsbqINN2qVPGgcf1kNI12+
bivZaBN1IB9WGZXiMQfJ0Pa6aaxiGAipxt1LtsGB9mfTZsoJLYxqeVZptT5cRziC
naAwdVKO5YwsVAygoJ0vqUcp6ePGri4s8M3LsXLyrv34jlPXP1vmrM/KfTdAgKBf
BI9Lbf/P22E0lz0N9mKgZRzmiWO03giio9knu6PV2Ip4Kx1WMyG3W2LFxvLiCElC
qOaS+Y/4nEr/hHFqmyHdmCwY5GJ8iWgTlvZgsn4z3xPtNcojH9/P2b039sMJgNHB
n3k9qd1myS2CEQVOF6frf41n+8nfrxXKk6k2YmtX6OOgX3eDQW6lqjUoEU+sQaV5
gd43AfxdDxycCJ6ebHLPm8UdMc+cXYF3eH22ctwEL4neIH4fAkzoeFZdMUxldZ0l
hbjo4uz/fALsHxoeyq60sFN2MfTArkEWhfAEyx93gigVhOBMgxfj6mzoKY8RJduG
ljetnuJoG2alKC2bRO9tgfEf2hUg7S+RQnPwxTNZynoV0PAyfsn4wnWMYw8WhN3T
yInuT/dP2SCMc/fqVuhlriMTg4KNAnN7BFhntoRKA+DXutu6r8tXldyzDLXJSCdU
QNFZe3ItCSuG4LVXtocjkV07mwKI4Gn4qVzrGMnu52lK6IkNJZANCrC13JPQUJlG
993hHUB27IiQ354nhYPt7O7vkY3Ke82ZKI1zg+c9AXB0uftXPYBwjRsuWMrf2b8S
30qpKOpR2I6SfSYKj/0pwuDOigHpVDQhaLdhhO+GH+0Tw+ZVyojElpML18fDI5QS
eUF2s574nODwuaK5mhQRJglR3L8+1/LzDsn2ITIeYxXgQ13cjvZ+7OYHjxfQKwp6
gs2SJItSZMChT5TQnlqTfA9kjVQ/fSAQ+q3oYx3wBK6D3j9s6af0/5iw1dZzx+ic
iouiek7Zjz4k64oVzGhUxtG8TFmDJD7qloPzkrcixWEFZLp95pcUVUWfJ5b6wQPo
cCnZelyEaQdTHa3K1xX2q6uRIYeC/KlzfKbItGlHoan3p/Y0ddhfSBJII5U1JDNn
uzCkRzROCE8s8d1B88k0eekh/nY8Omsd1oEtznDdYL02vz14ijxggQsiMFiCNAxg
rFx/iQF+PxHLhpzH95N0BWWKzGwaEeQYmzs/xGvBARdkWjbndjDpRgr66PKnvDru
kGw4uHaeQ+7uNmRatpu4WYhXiTHvjHumybPA2NGnip0jgkW5k7oABrZYKQBuAZaz
emxIM0FJSkW2/cameuGB5RDicpZEiR2cGszwUWDhy/D0BOFofQoTmwaYKpOaQgUi
Fj2ukYLLM6IW7v3KzB+B757SPBJUXTT0L4/cEacY9z68ELoZq+8xmNvziMG4TkAB
SvIIUN2lNibYzT9qZoh0a0CfS7eGwrLL34bPY3aWeIRYY1SZsa0FJ78jx1PNO+CN
m5n/mUH3UP9Kh/jsAojpprJsC+2iIrQdqzegH48fP80G7hZjgJP8dlf33qX18ySn
qJ2aWIr6OJuSMFOTgi/sHtJs2B3EW86rIYqq7hX3KHe+H91wPJ4GoZJDc6M6oosV
BgldF65x57Na5OfCx3C64sa7AJmAADgHpMG/3nCx1Z7eRnHozrOm4RQTUCDZiGKY
n7BeHnN5y6MgdGsTLmwI6vtPcPYSsFVLpe9ncnJtK3oUrnHbVx2xFMeZuu/7iMar
ufVFFmOPVmymyLbl0Xh5K8wLydU6i/Z5mvD6ZePQGxppe57K7hZx7euf8ZABzx6p
u26dZYnISRtawOO/sSsY48Ets3DkLZV1mtpPJNO7eN8SKe/KcnNTKuKMqAC/toNa
uIlkBGGPdVf9apchk3Utn3P7PEviS5MTgsrrNY9Agak5MfEteWjNbt70Z6vEoYz5
CMzK6G1zZR0thd3e3TTZmmpS93xgmChvVcT6lvb0lYTWxXDGaUxdsL6RmBUGGW4v
TcYfbVUh4JHPYByoJna6ZkprDmXEXQQPSnyVwhH4j1gv3bIbqPSfshgxbEKUIit6
Tz95WK5czl6eTquXGpEN6bSqCnswJPwNNwcn1aQyngqbshCaSC8wPOHzvkAtkNx0
lwYk3yciSFm/eTMxtqoe/kEdqX1K6fVqDQwQf/V9T0k1Dy5Hk+1rlXj1MQKFV1aj
n1+20kZdVO5RVmjNqgfeKtOaBswWfA1Hhc6d6pTpOxMkyLwdYdJj9VZtq+W+3c6Y
KNEt+V8czvSYsXdHuldpqNOAcn/kjrKM4nn4fP9cwId2P7Uqz173mqEOzaozopVj
LzRKxYSyf6BZLcZI+4MXIt8fRUxtO8BhC1GUpwPD4+CJgD5MQ5L2vuB75D3SNa2y
78ZR2mfSAaGIru4HaHtW1K+eqgXKExY6bKY9Z3B8OZdzr03abrF3Gnlk3fjkfddH
j9Orp1Tlf2idpy/yGEnRLcAJtwaRVzIXhuzfmbdQfVfuy7c/i4+6t78PE/SrjU+Q
geZVc/c3OBzbdXh/LX77l8DtnmJQhiNJnnXe/3QkWB3/u+jge5myRgNVTFdw9qRa
lLKgFSczsY3fbpl4D9A9GCbdD7CreAHvGn6wznXhmGLD7QUYMR3im20LiX54wZty
WzQ4TECym0yA68WvOIZUi1eT+w7pALoyuxIQWQrS3e5xDk/kFm0ky+guBWFM+Tfy
e25b0D3H6+3BQlToGfuvhsvBh2bfsMLzKxPKJ7mEpRPFTGKYAIwFAblS1y+kT336
i0u2xakwhoTXZsvgPdOYdFBoFH4RaMxlSaMA7ZFjVAK9Tu5SbQapkYYYsVwVwfOr
MSKfTyWSccfkfZSwMBBgHkmT/GWw9XLol0KBj9Z9vg+DwWxaMKlWfh/0tCz//jTg
gsQLmb5K+4my9L7LxYpffFlkTkWYkQRWzXGQlORK4q31qxGRppzod9e1sqjTvbkL
0nHzXCaa2jRXF1s8eXPkCK4lHzHTIT4XCW0EwUCDdORX8TCao0TriLxqyQfbpjEY
S7HXGMX5u81FmH8RfAlrt5mdh80c+st4g72yzh0koiZVKVL+GVV6khDnUmhmR5Z+
YQ8U0TKcoXDgV2XThzFarY95tt5d+aaUJZYvN46razrlT51gbzPvcBUfPNzo63k1
9o3TOk6ZmxZTvP4FQNT1b9+2CBlpSKkFxUORB5OyJ+MCfhQ+R5hEjVYtCr9yWctT
X36fipRoqpk4wDr1FENx6F1RM2pzLl9MLcnTFk1vEIgylHBAUsHKm3U+08/kk8Xm
lF6OuIKyCRhojuPuZqxQJ9/By+1zvXjlHyw/DrAIq8wPVJDEKo2+VeIyO5eh82db
LdbIVxmlR30vxuBCRLseKN8kL+oDvXd13OHY6NehDM/f2C6ZpzA7hVGgMxqJHAE5
cE1RcZOd4onKvda7ATawUxHyttux7dmIqLCGrZBQqNaaqENxJycboR2w5AhdwygZ
/jNM3ybKJTj/et+za+/Wo9UUAalXFJtcF+tfpSL9HzJekCfScsNdnIon3ylFBvWh
7oh7igCURPJyJvsoCLLjgYwbvcspBRNnuC0ce1gOaXLFPyJ9xZKnmzNQUakHsVow
lGenOUS8/zEOD4C+d4w/Q7m71HT4T2TJT72PmmTueXX5oQ5PdMNwPf01gkKF4pud
NIcjmBAs/7zpeXm0CBo/5B/EKApuhKQEmh/8GDHmS6r+HNqtteSq625RkwDwZnRI
2DYPlcF5MgnQRk9C6yAUxJSB1W/AJu3h2h/maRQHxjXCz3Lecs9D2y6uU7nb5S5k
LkBK0o59/FY89QM4KAo5oKpYS0RFmiyCr7aHL4UZy08QXBLCDT865Dw9zZrK6JQf
dRH8S0REGAordQKQlGQVvtDRSscQfspGVtI3gfx6EzYWmiXHuuvItFnnEUN65wcm
y88ERAEHQNYlqhERQ6fAm8PJ7/Lw1P73g5D+C2JXYdAeWNtRtE5WHRRf0CG7y5he
aBRaekAqkuwRM5qF9z4u/4WxewHK11X86OWGYVIbx0Z5sAXLOJ3Bq8VhA7A+9yAl
oGsiFoyFA7S/Kndk5JV5ZQVDTooGPxPRpSvy7huNKMwVaEffIwvWRXKVVcJt+7NE
rKbqRp2DSciNFRTMVP3Q9eyyPiwyLwiB6HRSWQYIIlysyW3zZSJOeuvmfqcKCsQm
65+Q07psQH9cSX3kCmYVY3RuW4T6tuVc9mhJakMdD02pAdL9V+W51NZcGvNoyIXY
Uk3xJaMLQYP0+KOOjAQZ+b5VcfSiizHI6GTmPdxoaMBwX8tRcJzxpAefE6fdlrth
c4IY+Cc/HE11P0F2v94PrvMO9uz2+aPSgVOODv2KSwKWUFrcNVt0YAEaabYuS7Yd
fPQbfJvcAcBY39fPGBEoONEeaRqsL1Kx2TlgXHH+s1VgZeCdn3sV6nQb39IxUs4n
j65xqvEgFMKy63awM73HCn/ShuYTAtisDRdA2sylp5VxJBTkEw8khzelZT5sUkEL
CwfBF016o6OEE70O/pjfHdMKqeAGBNL6ifV59Yb+5AuIj5ypjnWu9aJsojA8H+JB
jpVl/B3dJl3tCLEfGoH6OJM8OWPELOhCMO5MdjM1axoyEGdYztk4WbEj5CaPKgLG
2r+8kbeyH98K6bkQq7xXLAVB74KC5IPwB7CW+CfKthuFWMRlI6MEO0wQrm1eB16q
EV+Vn5XTvIiFqqC0i13FJc6jH678ph7so2A6A6VpyEM0poOKMvHHyk7Goo1xor6f
9QLDpFSB2mBR3LOq9gkBFhMu1AGFW0Vlaeikmxte2AhwsBSyhN9+K9FG6H/BSrVM
NcdKDJvMDME/fdyukt2l5p1v/E4U7QSzeCznxhEFp9zByhsaAPyIVSvKZZAO9SPz
sU3StGtX1YaKx42dpQ1AK/0h9DXzcy9YATBJIfvYqqlQ8pA5N7VYNqx8AoOWkTYz
noaz1jX6ots7RrxhHRknsRHewYyAB0TWDEF7usCtyYFBDq3885AK/oX/hB5U7VeQ
Yrt8poc0cY7O+Hu8VM5c1Txz9bwK3ITWOfD/QkBZdPZ3USEg6KOP5TIgqJW7D+RM
2/kJZyKHfQ80mGyYgsG6fF6ClamSpo0ksoQns9lcdSs97CXT+6F8vvPO4dvS90fu
iNP6f1tQcXNhCEugSrKe0Uk8KHaIyYC57vPg7sMsUh+1W5OU71HN03tyz/WV+T/N
RnfTkt3C5ox+Za7chLU8H3HFKztKH4gOsl8r+hnWi2wkiukhlo6nyji0rXG8GdOz
6F/3SDhI1yZz0ybdwkzIRofCRLJny6c8pA9JP/JBvxulbCietqr0q5ERLuYfo7qR
4Ki+Lqb/oxyeQj1/bqErw7PhTy2vToVdCc3x1BkpQQGPpFEQ51HBEgjefKhg8p41
1tkVDAz9GFNIGJp56h87iG7CqpXw8IOcb3oxsBq/K1FS5XI1kkAa8N21jZl0fayT
OpknS4TiOu/kg/lPTMHl9XHI7DEgrGQMriHvPwJx+TkVIjEZB0KwfM7SWaB13kQP
is/uW8iNeg62Qith/ad1ouonUoBO8ZvpQFKRjlMhBOWYsYKze7hS2fBwmi3WdKkt
B29s7dVPBqKO63tYC+GW4J7MrI0CUziNq2Xgr6TQiDM0RTUIZx6vpfD4qeGLss1Z
0mbiCp8NUQtaxYtVZx5rCr9srHpo/XeCy4uJJQ3JGW5P1xbanwL4xdgL6UCo8qhg
7eoIm2ycSTGfq1F/2PKA3iCikpgSVgkG7Zsu4xwWslUmBKUSabgnDdXwEEhZA+Tx
1rx2IxPhwJQ6EXBkPrL5jODxO15uWwCYISuYIlzwJxlQZhgST/BgrzVVL1Zi+Rua
FYbj/AjizxXr2Nw24v3v3nNfUt70QXMBZL7IrB+bd0Ukh+qdZRdDBSGwAZAUCYIH
kvJweKKE8q59DbPvgRggQ+ZRwkQsQWOxjjE/GQMOxonztHoIA60VZkpZfXfQ86/s
yClmzMCDknYH6GIYXvlPV0KNT2Umr0nQw6lyMxkZZIGMQLkJFwdmZt/PgIXQrMGB
2cQsS74LLy4/cN23HqiuG/TldzsVYj13f3WKp8XV1qB3lyflvi6IdcilUd37avze
m2FDpkJLgdXYe3Vu1a15fNmM93Mh8JlvJfMD9nxNf8DhaJzMFcGX/2nmL6mnonJs
z2+97+y4vtL/ozQatzjAXVdd0V6DQ5WlQkKt9mh5Vwa2aONoFqscOK/0oP9Q1wUx
0s+rGdjMwimzGf/GP5cPU0caXNnVz+8dKSwsjRyk7szm0+B6qRJX1QiXOqNyeQkA
Z9QG2/Ja5Mfo5aTiNdX+rDU/fUd8Of+iSHgNpfSjHdhrDxVZs9k166JmFcHzrvZ3
6ACRfrjGlLW5k3Z4z8xQ9XVs29y9YW2V1w79n7UL5ux7ICh2KSI2Xw5deCDs2/9q
S9BUTtnl85jfPGNFMAbcJ+FXUntk8oYmetFVFV72v3lgm4vJt2GjQJwqwcHp5der
0WEMkfNgiZre6QoFval79I2ApzlXsnx08AT7tBOIl3NxoWxV4FiwlgbVVQLfM9tc
z56WU3Q6nEGi9tYztlRIUY4pLTNTHc1OJfBwafUgp8BojXvxczpgOzwdQw2vVrCv
9WkLDTj+ho/2yld673gBKOOPZG0ftJFU0M5k+gs17lpYt0OucLDmqwxY/jOe0RNJ
sqPFMPFOT4cnYunLaYO0lSCyy/fcBM6hBFQkr3BMQFMFdN6Wor5zqfaaurP4o3lT
H6sKltsveWQ/jLjaAmlih6GcauX1I6tnPBGbPla5Di9IGm5u/fIkjya7waY82MMc
1+JSsuOHYIjSCbQ1tHgsp00lSV2FOineC/oMSnLLJDHZHN6jfdmlJ6mDHnFVXVEn
C4jgIRTuKuLFuFKmAdCi3R7ccftS533yvZv6dCWFQ9ie5B5YlgFau+h+pjvKgsEP
Zk9qcLA1KCCYQK6WwM62zMurjAbASeNKN2dEw1NYE83Rq5F2iGcewgdg3wgDEgze
wmyK0h97YhZ9f87xn7BU/PXivRD+gE/+8QSkRfvRpgN6eVR09VSjwmWjKH+1Qjgu
5G58nUAb6bsWMFmeEqLIeT0/uqfKixYKBMMjtj0YmchnCIZw37Qh82Jwac3R+ETP
VHJLRmKkdjOb2+MGB8kSvMzulv4zb6Nyf/b2I/7Mu1FnN+cK4uHqSYfL7vlIxDjL
CA536TY9aEOteSm4vIBDHYAyqYMDDNbZ6gXtUOUmH+nHNzWZEBYcypoNbxr3QDeY
lKM5CdjZJIkWlfJbxqQVw6oloKPYutjzg2FMTz5AA0WDAJ6IaPxIsN9Mn8CkIDBI
SkSfixsVacwDI6X87QwNNJkBqqH3bwArgBakzZ/9tNxspY7quJzcAZHKLgy1s/3Q
xJrTqgt9JqQoX8NB8VwuJXfqo826CLN7jW/s8epysje58Uuql6IpEjjyM/RDr9ts
qpp1Kz2fjhploLdHAE+agTEbZNcVgP7zyrqsd8LIUvgo53pT2jukc6VFbMPqqVW6
K19eykkYeinBSgY4GJZ7kw==
`pragma protect end_protected
