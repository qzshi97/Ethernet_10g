// megafunction wizard: %Ethernet 10G MAC v17.1%
// GENERATION: XML
// Eth_10gmac.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module Eth_10gmac (
		input  wire        csr_clk_clk,                     //                    csr_clk.clk
		input  wire        csr_reset_reset_n,               //                  csr_reset.reset_n
		input  wire [12:0] csr_address,                     //                        csr.address
		output wire        csr_waitrequest,                 //                           .waitrequest
		input  wire        csr_read,                        //                           .read
		output wire [31:0] csr_readdata,                    //                           .readdata
		input  wire        csr_write,                       //                           .write
		input  wire [31:0] csr_writedata,                   //                           .writedata
		input  wire        tx_clk_clk,                      //                     tx_clk.clk
		input  wire        tx_reset_reset_n,                //                   tx_reset.reset_n
		input  wire        avalon_st_tx_startofpacket,      //               avalon_st_tx.startofpacket
		input  wire        avalon_st_tx_valid,              //                           .valid
		input  wire [63:0] avalon_st_tx_data,               //                           .data
		input  wire [2:0]  avalon_st_tx_empty,              //                           .empty
		output wire        avalon_st_tx_ready,              //                           .ready
		input  wire [0:0]  avalon_st_tx_error,              //                           .error
		input  wire        avalon_st_tx_endofpacket,        //                           .endofpacket
		input  wire [1:0]  avalon_st_pause_data,            //            avalon_st_pause.data
		output wire [71:0] xgmii_tx_data,                   //                   xgmii_tx.data
		input  wire        rx_clk_clk,                      //                     rx_clk.clk
		input  wire        rx_reset_reset_n,                //                   rx_reset.reset_n
		input  wire [71:0] xgmii_rx_data,                   //                   xgmii_rx.data
		output wire        avalon_st_rx_startofpacket,      //               avalon_st_rx.startofpacket
		output wire        avalon_st_rx_endofpacket,        //                           .endofpacket
		output wire        avalon_st_rx_valid,              //                           .valid
		input  wire        avalon_st_rx_ready,              //                           .ready
		output wire [63:0] avalon_st_rx_data,               //                           .data
		output wire [2:0]  avalon_st_rx_empty,              //                           .empty
		output wire [5:0]  avalon_st_rx_error,              //                           .error
		output wire        avalon_st_rxstatus_valid,        //         avalon_st_rxstatus.valid
		output wire [39:0] avalon_st_rxstatus_data,         //                           .data
		output wire [6:0]  avalon_st_rxstatus_error,        //                           .error
		output wire [1:0]  link_fault_status_xgmii_rx_data  // link_fault_status_xgmii_rx.data
	);

	Eth_10gmac_0002 eth_10gmac_inst (
		.csr_clk_clk                     (csr_clk_clk),                     //                    csr_clk.clk
		.csr_reset_reset_n               (csr_reset_reset_n),               //                  csr_reset.reset_n
		.csr_address                     (csr_address),                     //                        csr.address
		.csr_waitrequest                 (csr_waitrequest),                 //                           .waitrequest
		.csr_read                        (csr_read),                        //                           .read
		.csr_readdata                    (csr_readdata),                    //                           .readdata
		.csr_write                       (csr_write),                       //                           .write
		.csr_writedata                   (csr_writedata),                   //                           .writedata
		.tx_clk_clk                      (tx_clk_clk),                      //                     tx_clk.clk
		.tx_reset_reset_n                (tx_reset_reset_n),                //                   tx_reset.reset_n
		.avalon_st_tx_startofpacket      (avalon_st_tx_startofpacket),      //               avalon_st_tx.startofpacket
		.avalon_st_tx_valid              (avalon_st_tx_valid),              //                           .valid
		.avalon_st_tx_data               (avalon_st_tx_data),               //                           .data
		.avalon_st_tx_empty              (avalon_st_tx_empty),              //                           .empty
		.avalon_st_tx_ready              (avalon_st_tx_ready),              //                           .ready
		.avalon_st_tx_error              (avalon_st_tx_error),              //                           .error
		.avalon_st_tx_endofpacket        (avalon_st_tx_endofpacket),        //                           .endofpacket
		.avalon_st_pause_data            (avalon_st_pause_data),            //            avalon_st_pause.data
		.xgmii_tx_data                   (xgmii_tx_data),                   //                   xgmii_tx.data
		.rx_clk_clk                      (rx_clk_clk),                      //                     rx_clk.clk
		.rx_reset_reset_n                (rx_reset_reset_n),                //                   rx_reset.reset_n
		.xgmii_rx_data                   (xgmii_rx_data),                   //                   xgmii_rx.data
		.avalon_st_rx_startofpacket      (avalon_st_rx_startofpacket),      //               avalon_st_rx.startofpacket
		.avalon_st_rx_endofpacket        (avalon_st_rx_endofpacket),        //                           .endofpacket
		.avalon_st_rx_valid              (avalon_st_rx_valid),              //                           .valid
		.avalon_st_rx_ready              (avalon_st_rx_ready),              //                           .ready
		.avalon_st_rx_data               (avalon_st_rx_data),               //                           .data
		.avalon_st_rx_empty              (avalon_st_rx_empty),              //                           .empty
		.avalon_st_rx_error              (avalon_st_rx_error),              //                           .error
		.avalon_st_rxstatus_valid        (avalon_st_rxstatus_valid),        //         avalon_st_rxstatus.valid
		.avalon_st_rxstatus_data         (avalon_st_rxstatus_data),         //                           .data
		.avalon_st_rxstatus_error        (avalon_st_rxstatus_error),        //                           .error
		.link_fault_status_xgmii_rx_data (link_fault_status_xgmii_rx_data)  // link_fault_status_xgmii_rx.data
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_eth_10g_mac" version="17.1" >
// Retrieval info: 	<generic name="DEVICE_FAMILY" value="Stratix V" />
// Retrieval info: 	<generic name="ENABLE_TIMESTAMPING" value="0" />
// Retrieval info: 	<generic name="ENABLE_PTP_1STEP" value="0" />
// Retrieval info: 	<generic name="TSTAMP_FP_WIDTH" value="4" />
// Retrieval info: 	<generic name="PREAMBLE_PASSTHROUGH" value="0" />
// Retrieval info: 	<generic name="ENABLE_PFC" value="0" />
// Retrieval info: 	<generic name="PFC_PRIORITY_NUM" value="8" />
// Retrieval info: 	<generic name="DATAPATH_OPTION" value="3" />
// Retrieval info: 	<generic name="ENABLE_SUPP_ADDR" value="0" />
// Retrieval info: 	<generic name="INSTANTIATE_TX_CRC" value="1" />
// Retrieval info: 	<generic name="INSTANTIATE_STATISTICS" value="0" />
// Retrieval info: 	<generic name="REGISTER_BASED_STATISTICS" value="0" />
// Retrieval info: 	<generic name="ENABLE_1G10G_MAC" value="0" />
// Retrieval info: 	<generic name="ENABLE_UNIDIRECTIONAL" value="0" />
// Retrieval info: 	<generic name="AUTO_DEVICE" value="5SEE9F45C2" />
// Retrieval info: 	<generic name="AUTO_DEVICE_SPEEDGRADE" value="2_H2" />
// Retrieval info: </instance>
// IPFS_FILES : Eth_10gmac.vo
// RELATED_FILES: Eth_10gmac.v, Eth_10gmac_0002.v, altera_merlin_master_translator.sv, altera_avalon_mm_bridge.v, altera_eth_default_slave.v, altera_eth_10g_tx_register_map.v, altera_avalon_st_clock_crosser.v, altera_eth_packet_underflow_control.v, altera_eth_pad_inserter.v, altera_eth_pkt_backpressure_control.v, altera_eth_pause_beat_conversion.v, altera_eth_pause_controller.v, altera_eth_pause_ctrl_gen.v, altera_eth_pause_gen.v, Eth_10gmac_tx_st_pause_ctrl_error_adapter.sv, Eth_10gmac_tx_st_mux_flow_control_user_frame.sv, altera_eth_address_inserter.v, altera_eth_crc.v, crc32.v, gf_mult32_kc.v, altera_avalon_st_pipeline_stage.sv, altera_avalon_st_pipeline_base.v, altera_eth_packet_formatter.v, altera_eth_xgmii_termination.v, Eth_10gmac_tx_st_timing_adapter_splitter_in.sv, altera_avalon_st_splitter.sv, Eth_10gmac_tx_st_timing_adapter_splitter_out_0.sv, altera_eth_link_fault_generation.v, altera_eth_10g_rx_register_map.v, altera_eth_link_fault_detection.v, altera_eth_lane_decoder.v, Eth_10gmac_rx_st_timing_adapter_frame_status_in.sv, altera_eth_frame_decoder.v, altera_eth_frame_decoder_pipeline_stage.sv, altera_eth_frame_decoder_pipeline_base.v, Eth_10gmac_rx_timing_adapter_frame_status_out_frame_decoder.sv, altera_eth_frame_status_merger.v, altera_eth_crc_pad_rem.v, altera_eth_crc_rem.v, altera_packet_stripper.v, altera_eth_crc_pad_rem_pipeline_stage.sv, altera_eth_crc_pad_rem_pipeline_base.v, altera_eth_packet_overflow_control.v, altera_avalon_st_delay.sv, Eth_10gmac_rx_st_error_adapter_stat.sv, Eth_10gmac_txrx_timing_adapter_link_fault_status_rx.sv, Eth_10gmac_txrx_timing_adapter_link_fault_status_export.sv, altera_avalon_dc_fifo.v, altera_dcfifo_synchronizer_bundle.v, altera_std_synchronizer_nocut.v, Eth_10gmac_rxtx_timing_adapter_pauselen_rx.sv, Eth_10gmac_rxtx_timing_adapter_pauselen_tx.sv, Eth_10gmac_mm_interconnect_0.v, Eth_10gmac_mm_interconnect_1.v, Eth_10gmac_mm_interconnect_2.v, altera_reset_controller.v, altera_reset_synchronizer.v, altera_merlin_slave_translator.sv, altera_merlin_master_agent.sv, altera_merlin_slave_agent.sv, altera_merlin_burst_uncompressor.sv, altera_avalon_sc_fifo.v, Eth_10gmac_mm_interconnect_0_router.sv, Eth_10gmac_mm_interconnect_0_router_001.sv, altera_merlin_traffic_limiter.sv, altera_merlin_reorder_memory.sv, Eth_10gmac_mm_interconnect_0_cmd_demux.sv, Eth_10gmac_mm_interconnect_0_cmd_mux.sv, altera_merlin_arbitrator.sv, Eth_10gmac_mm_interconnect_0_rsp_demux.sv, Eth_10gmac_mm_interconnect_0_rsp_mux.sv, altera_avalon_st_handshake_clock_crosser.v, Eth_10gmac_mm_interconnect_0_avalon_st_adapter.v, Eth_10gmac_mm_interconnect_1_router.sv, Eth_10gmac_mm_interconnect_1_router_001.sv, Eth_10gmac_mm_interconnect_1_cmd_demux.sv, Eth_10gmac_mm_interconnect_1_cmd_mux.sv, Eth_10gmac_mm_interconnect_1_rsp_demux.sv, Eth_10gmac_mm_interconnect_1_rsp_mux.sv, Eth_10gmac_mm_interconnect_2_router.sv, Eth_10gmac_mm_interconnect_0_avalon_st_adapter_error_adapter_0.sv
