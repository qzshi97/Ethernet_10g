// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:28:49 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l4HGhlRH9wWET1OEXyibgaqYKtx1jR+y2i5qRUmZ1YvxF7rwzwwBcjVq04k3614E
utpTC8AHDZuB3POr7Ua5+WxCSAGlwAOVQdvaFChT59t3ZfBsU7dA4cN9EXjQpDYk
Lfy5OHGP166tez9N2HmkCnCXfVRJ7neUNdQqNecTl1E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22672)
qWq3QztO0ZOwzy4I8dCD7ODQGIqEaOwwmg6F13ypI3okstpVS6S9x6YJ7w75JVeh
NYdMOkuFEts0X/LSe96Er9EHhnde1kPIr8KxDXtQJ6T5CpRc76fEDx9G+vK4LWcW
CT2502gPwXt2rr5qxnp41ImcASF2HLTAti2ros0WuDO0y8CAtdqYudS6DI5Tsaw3
RZZN507lD8ivug39mbpJWr9zCzlK/uGD6bQu1uAm2NkfUIIJc1l9iTtr4UWBWNLc
EyjV700QwHnuQB6mMUZhoviZcL2KVabpGc+EJTrCuSj0JQF+LqoibnV1ZzKbFGMf
lqQRffa00qawXZoUGl4nq8CdEfLqsxvorki4x0tjbsOSBPnxcp5ZEyeuGLq8XhvT
O5PlPejLWHzH4+xEGUu6CDgc8uXkyR107POfu7JsP2iciPJhXwdVT2/Md51aGAV/
pGNNqMCSF1DjJIXu0IcQKTsn90DOAyxPeNNZv7p/uYH85bmDas83jRrzfBYvjP95
pCKljns9rB4f/JKAW+SiDfJl2Uu+9qJFIfObiiJFGTRrqf2gw5/XTGThLaabElR5
KSC6BwmAc6U6XCU890yR+l6AaiTPSXazEZxy59FyjgciSJKjjWMxVufILJQf2x8F
mV9id72HQly4WT9PJjS5Vkfr2MsLWkhMztvWjMcNEnS/Zoh0k7fzt4LN79iXV1PB
sANXEHp63Wn3pQfc//ckiBnWLqk3D3BtmTBRxryTJgmQpiyKPkDejzYxvzsftLxs
/McvMFi+1XoDzEEG2UZoEFN4zN1Esl5vTOJ28vWNF5ND6Nek7FzLumzrHMCUXXBd
fSR3IZGX7gRDkICQlvqRygphNem2bV2paLYT/h29p/4ydXJzA614AhJwWZ+LN62j
J+fq9O/P+2bkl2eVfpaXvaVZ6Yx11uGbDtGOvf5ZtpbmO8stExT+dhFUJqYvBfrr
N4WlwHenpLw2zHnVj6jkszAnHjLmAc2E3QaVX6B5QOGefL3RpEZNk+zcI+nYiN5m
uIq6jHFTNoR1vyZ5m51jChTI8LDzplhIQgDoeq4ufzIGZ/wt/oxBWZqyyDWVcUIW
DQU5zZ3VBmLgOcCQOTcdA0aa3AoXidv/kMGxeKaFlwlxnmQemabP0OKy9ihODGez
0p4tamBt+zDbaJ7NPncMzTV3AZLP4L5pAbAPAhM0rcW+vPBIQ+4GfNcdBXhRVa0u
dx7VHoycTIPsNBHLSlmoVzD9CSQXr70KcjGV0aYCn6GAEwhwMZ/vwKkQF9tAfj1L
tl+MV7fNeKxW0EOnO1j5YAdfs4YxN3m3cZBehk1ErdeBMdqGs89Prrn0IDoEK5UR
ZLfCQRp/vlYyYKzERFferjMMMhAdK081yLnj185R5uDWs8/kaXQZ2wmd/u6jdeNB
hDp42NPuG88ry4RtI3bJlmGmzPCnRI8FJQiwPp7BKgWmmWg3f20p8qutT/7+WSYk
DLIfhGOB2bEquPZ2upIBziJBSKTCvS5v/AmkEjiLhj/NA7a95e0VhkPk22fieUdl
bvjhOEKBdwB/Io6r4McLA+5LOo/2xc/WA7/y5g7uTLv59vfTSb190TrTZvo8M93o
wGjwb668Kq1qJ36e+pSclqD4H+cNARK3o+bqXnLcJh32eGsD99ZutUlrvyEBb7DH
FMk7gyFZiXOMSWkK9/HBNKs7XD7VN8mjoHnkSsaZpiycRjeStRQVr0JKxIizk0Ap
f3omu9RdjsuZ0kT6EzDE0ZZpkXOSYVTUygokOVYxdTx1YmAlrEHvYuZYxpcxdFKD
Ih+T2G+R7YyinVnPy3fXDnz9ch74TvMjQymxwaPWRUzGjuDBI7nUKr0dhkoxNcis
IG31WUsBfIKfzaIcycZ6APiK5rAgb4T907XAmFKUjXWkHbreUBhsmUyXcvv4VKAb
oRr6bjD64qEECLoppQy1o4NMdF/ghEnFalihRwYQI19a2HxlALg8ciRcMv3L/KsZ
1v5Kqggh5H7DAsvs8hPnhAVC6BuD2FSanQWty8rjd7sVIPN27vXyOz/Ed2H2zEab
lGzCYKQPMWn3h2PuskYcpCli75mVc/D9adeo95tBASyI3Xz+8gKJEWvAk+27xsp/
BwEysN9eHfaoTV2k2NnOf+NgJvP9d3pcHZwWnmiO3OA+fF5NymYJ4FU7KzUZg4oE
4HlF21o3ZLT3J6tjmFw3/CN1leExZN7X3S2cw/rxCWFRebjthe8ZTKMsDibq8jNa
z1JMZjMk2C52zLm/0YOEnUFNFwbrB6jKbHAwvFsmYJsT2cCcjUO7RRlt20ZimP5O
y8GhRhqZLX707CTJWHwGRa7t/ZkCwpM0qybfv9e+p2bcidMHwhG6cTDL8j71QmeU
o4n3Y/ESf4MCPMJlcr6MrJv4QPvLjSsZl8D9YELTJ+Bu4eQSVJKu4NSkhX/EwIdy
USEVhFedVyrrpUYwTYuBjrS2qYm7y+K+FloklFndNhoUzHINkVNbVA9mOiYTNz9n
A8HprJsBB0rjq7DHddHKavpogPIyJXVXtpHYZzzKRt3NvH6acWdTAZQpCfJxepvI
j3fwjenJ2/8Wqd+ucnLeuIujzsjYyUf7S1uS/DuRIiQqhSOZtZK/M5C0u0USOBuu
1gfdCCUVGQT1bOtan/41pYBvQk8zpQ/T4CDibU1mV2A1aGixPmvUIoR1tSEj+uVn
bBQzrtRMBGYh1BJbu7iHZa+Z7AsvqgTYhnjvlNU2VZY8xt81NQFsEydTXKHJH6nK
FufbUa2cyXI/BYgNedo7AZ8E1UUXQYcDEkbresj6ZsLHNMeinmiYfo0s9mCNV2nw
I08JP5Qbo9baS77msg6m5hoUNUEScfVFQyfr6cAoWfFdPJ/4A9ltOxMs6dSCQIP0
uON4oVL6OuPG0Gldt1UcB2MXaIZ4zo9S1zIvmBdfCCacEmNuRe68SyuhjKdle2Sb
Pl2qBl001gVFNYyq1/nrEK3kQu793LB1zSKtMpMCMtQtU7Bcw4RZ+ErnH3x88o54
2D5mhP3bndXnNJHrGNU8ReVrRV0JRGD4oabRTKgIOw/xm+W5N+/xCdjMzhCmWhhx
obX5fJz7GnEYfhINoJVU0BPmwyLZWaiU62YkWNzmI4Wn4tXPveAs4SCt3iJalGG9
gjlgx5af4bvLimH0JiVUcaSwH+KCMLr614S0Oas10HYlXDzaTld+LCooshOj4vlT
V7iS4iHqBj1rHhL8NyBLbRe7sveL09wpyVURsfvpDjK84RX/XzaFAVs0uawIdf6g
cUS9NvMKGQF1MHLUEv/VC4cDbKKPRvtRun82O7gF6QBu4ToAI1BR3iuww9Mcmsk4
A8MYAK2HyGSB+rHfoItePa9fUFbuNlaV4JzrpF84wSMAbUp4pJxIMcJrLCB9KUDY
d/K+EBx5fKYvSvmIPS+aBs6WfpvFUJSoxpSdbU+6K8r17shx0yZyB/qAq2jLIBXy
gYuceCrJSxMXXoinU7aCwTKfjDuE3zrx+/Z8owC8ImxP0A/gAraQCi1fHrslFqsL
eZsHyu9Ex7Nux7Fc3WrZRsCZugRLk4c3Wk2mHHiMomjs27XxjiQpKXuPTi76fgz8
hDj3HHfOImtxojO2mz0xTCQAfy9OnPaY92aa09OIISy9SO6+vtf4aJlP5hSUcBD3
kZYojeMHQ+yYt3ZxNGQohQM6khtHkU6ouStOFdXyS2kO0EzbvZL6tfwA2heQDC16
Xyq7gSiJr0caEkrmkuA1r8sv/kwk0YySv+sE63n/D50AY8XRbLOQwJy5MPOtZhFh
hdO+No1GTRbJVTqMU2ODzAA/U8872FKmi38IFVceu0/wrW3aphboOadrnBHdbTSS
XnVVcbyppeCg1MO7Ct3WFbqVQEEOt+Z96blQ8WCrD59RGkO3KP26GccWQfa2SHaa
1leaoDPY/gQsnAXjMhCJ7SHcZ3qYghgmvMzUEkzMCiyTvHPOqBAoE8Rd2Xgkneq7
c+DMncvPJdOVhbK0Gk4yZ9HCeH5GWlFaW0WWZHQwUFyUysHMm7pdl/gF0qF4h1mT
ChmzJAPaIoUOeDnoRLx7hrNqPKuop/F4NrnU7i/+YGixLIpulBLGOwlZkrj/o+h9
lH1ZJaP2dsncE3xcEJDwfAqIAZNE9YRjth/XhT79tX8ejJ9d0JcmLehD9zB+vpCC
41xgp8u20/BOugVjTOzBZAqgHSK/0ujTJxWgu2ORfYWW/XUBCTg36wM+PwUMioPZ
+8zxC6N+8zVGh2IAUYQThtEl4u1p4piOP9AbL4LIDtzH0wIEDEfnlGoN5ipOqpDt
kaM0PnuP7ODfaFyRGpPc24+qNAsj5LUMLfXyer0XBkcS6Gs7FZebxZMdyFqGC10U
Vca0ZmfNWK0CQ5mVKwWWWZIjyjRE9jaLUe4Lq64cnoGJ62zfDm3Thj0JuTTqY2hI
YpuyiNh1b592SmlV6Ym5sXO8eZG8bsNBRCx3/sQQ8Pf21nDFop5/M2uxqg3XP3YD
W0I25H3IXj/Nt3/9mf7UdjBxZtJw15mZfdb4JW5d21EV0WY9njUu0PESXbf/5WDd
c4y6U1YMSSUf7ra1MygiM/p9L7OCiEbQxaqO22NZsNI0YOECNzaE1asYvgC9hh6A
9dw4Z+7uoiQWRAaubpm4kZfjkew0BpgYH+PpCccvoLFlmdqc8MCh+v0fRN2b64u8
yx0nzE/7fMGoE6Eyi8PuGDfh2W4aBq1GF9iWulssa/1qwjwrj7xg9q6xm9vnQAkl
uFAYeOT03OaT88LMkpCtszRmNVggw39x/nn4GY/DznGbJCpbprMHGGhqPHYwHIw+
nAxYq1VkRXTeuOZjLZzN0ytplTLl4wVLK0ZOgkem/RsYU5ElpY9FONBMZKmmoTDg
d48tuvUKwBEVaHynsmqlT+s8Azr3/uuo0dV1GMVc4naxsuZPCSiBywSHtk8xqkPI
XYUxspY2B9iol0NUqWwxPPhQOvi+yM97rlyztw2vxCoz5IRdAnUgtkIvzeMPJaf+
18ojR1gsPb4harM9qWruXwu/iEpT2/sBIJKHrjNvA3ruB2ZYG/6Z4Nd5V2fY+uox
Kk7RomPJKj6L6TGyUOnlmuN2+AWQhYf537vJn1oqywFUz4eACFKW1E+wszuDElLh
uVa4LgUpvo0SL8/5q6ks4JrIH0YByXkl19HKr8ul8rnzqe7QUBOgYnlHJ1406MC3
hmvciJukBS3NJeQZm6PFhsArQKRfyxWYeyR+uFZccnTlvixbRAgImER3j3va9u2Y
ZoVUvA9X0gXAvk6dpMyoZMbkpf4UAz+kC8kJlBU8VSk10LLVRPaM+/EpqCJ+3T1R
3GEuF3M7KUoWby4wfrZweRk5b/cz2L2wu2gY8t14dqrROBY8R7z+OuEo7VoKyTC2
U1nOK5iMf7ta4zD9BOPlI2NDM5/8AiB/5LiJerdTybKYsaoMxFyVLFKnLbLwW/Fk
sUq3hZ7AftxIag2EPkYyn7T57hMoJYea50j7P0W/88SLoJxrYYFfXYwa1bIYvUuV
wSlRJ6ZrKtt8leIODSQFAD814k3ktgRhdx1hf5r6GQR6uxWRsunF3Hgk83S1zu50
iW/lXLeNP1BiPtQy2ywYeCje03FVD4cgF/wut9mmYvaOXJ2iZCSMa+3UDg6e5EYm
M5vQt2cGXbOewSH6MUREqlZkxtT0AKTMqZ0Hkh5ZNe8nio3fKBDnKoTtkzxuOvoX
DrVhEA3NEwMlsApEZdnWjHEAAf0OdhFrj+iwP1S8sAmIvH+V1oepjxNK3yDPRfW3
Pox/JTcLWTfBO9B5ixDkzGu3EOfKVwAIeHCYNt+7WcFNUOaNz7FNRk4NFGmTJKqS
TrKwnAXUfC2o4NZREKnLwL5qUBPJmoecQK4CK16E/KalKZq+DKMd6r6/Qul6LJOW
2KXOOevo6wbnWj383iUeXP/m4hwQHMdhYUgJv3OLPiPwTG/ZDnMWPB79SZgoJC6s
Gwh/HGl9g5yW/ZBe0anOTNq9J5V+4eZlMAosI4JqkspSM18Un+dLEMA9gR4bGpFl
KCuclugR48xRZpoc0M/OJgeq23t4JHpZdqxUUqRgCoD6fLL6F4UrgX032ylAq+gI
ScRx12tmKybW5/5csOcgoPqXcJEdsU1u+pGQaUn7W+FYakii1y2UGGQF9qo0uzOF
fWk3SsyOTmWNPxbeeV3to4rcOZcNGfudWbMDLAWapOmIibqUjGWGlHBFrhnlwQj2
NiCJMFQFdKmDF7wCkaGoySHyGsJbFuDF7UcU6HPRid5jOK6DTC58dPixqY/mgJ2L
Crvye35E6eEFDN/BhOp+XVgkykwIycYej3NDoE1oZloQbja3wD7hEQOFGe3vtVjh
I8ANHK5msR6iRXRbanxGQ77PQNhaiFIiRgusciB0Vc1SAaT0nucOQY+mXMUjB9sD
ntojPuN1cunHgX8UpwhuYxFm3T46qnSNtu09rSCfsNfwpuXHSOVcxwcjm+8sr+om
+8Gp6bMW7Ij51kbFXPi5E7WY30RLV4YgHDArpwDCEOMVIrz2Q+6V78WkG7IqDi70
EEbN08otxM6zdjRodyP1/BwVCahhdIfWlNn9q6iQFWTPdc9OaLzPA8e6N4dHgipx
cCFjLhIWWNVZvkRU5p6VXcJV9JoyJ9kMQFPKM0aFld5MiGUvqNG6E9fAk+B444fP
UxQXBG1jYvg5RixqUFnwLBC6XVnpXrzvHccNCjUYmxxRk2v2I1n8pebDJONk5uJm
0p/8dTfoCFVIJRctDQhdSei2kwoKqEXDE9udmclZdoTxkYHaBwn06Mgs2OasCh08
4EDTEAwm71DV/Nno8PXyi7d8JrltA2uyVDtIizYgW5FG1r/Pvj9GY0Hvb302aJkO
UU9ks6Ei82OR+oTzHo1e6UiqW8GwXH5tbDvblIXEOfBdWkSUPqFjdTLKy7VpxtoJ
KaRdU9w1ndlwv/ceEoqwxzGgd+y0RwtRzkOwA+PUjRuUPxLus+1UXX/TgZjoZClR
2goxA6mf/GJMKlRvUVQZ9zzvADWGDyXiacuqBwG7RQWxjrsSUvDo3cVz06Sc8CyQ
0JY9wckMnfwQ9G/mHecJwNBti658NEYnzvqgzsZT4yYPMglv3vBYzgQEkEI66PW8
6Co/Zd8ReyCdco4aDp6yey2XZPuy03VLIk+JvVg0WXB75Hs3XcOQU/gLsXdHt8gy
fGqArPVAw3pMkIDiD+YBobw95D+MM4EUNtapQ2E1UCre9d/TAi+iBmzWL8OK49Fh
EfrrpGivaoJG43yJNvs1GewCTB8/SD8MAfv3mH13JCbZNPhL7YSjqLqesd2cHYiK
JAK+bPhTy0HovtGqw4jspCtP5qdLGU8IyErNiCXCcNLgxO9qHYCWzmCeHPuWsOzg
tzAAQKwq4j6bR4mF1sfeZ3A+9OW0CSJItuY7WVnUo9fcQZ7FQ4KHXOC2FbWNiKWV
KZepA86DhYpAysfEKfCEAM3TWzQaDT7aU2AjmI8gMMfgiBsVRbQdH4z56vT0Xym0
WV+G3TUJjrwMTn7lAIXbRUZx+JOIN0saiL9frk29bYlzVZot2KfDMBhuIUhdxR/8
1s/b9EyGVgRH1z62hUqFJWoHsrE47Q9Ta7140vMESYmXHeJ/za7sKpmW2SfLD9OE
pS76fHISW4vxVoGGzUo6z9VxfULs9wElc9U3G8SFpWIBi5iv8cTK/kCtU2PB3UL1
s+2YNerW7EgZZZ1Lj2nM0Z4M4zYgceSJdcn2LAFALsyS/eD7aZm5wUYVqZHuK0Ci
DUMY99zSUOFZqnm/L9CsrvKzvlnranOIwZexwOPn9NPuookWe4CRUDNXmf+GlixW
tLJClEYUUJVL2FxCLg51qHqeF4YwNDSl3tfqwCCYfV0kngp1rUzOv5At1Q6ie5vi
FZ6HFzRuGisKsc43B9RUbzBfM6bJ4d57xfTLNN/2PGzPu1Pt4BF6yVoxvDkA4CHS
KeEvUtdZEpDaoxNOfkDK/eD/nml00GqJwmK69H+y6k41YjQwDiFL5JlDoYZMjl4R
F8rsAmaOjGGJmKGc/sidBjQO+bjIYADRtshEiDQES9pq/A6fHlNKV9qL7ubH/0h+
uktO+N8SXPZz1H91NuUHUkWhqdL3dm5KQQ9feilh75E7m2aP+9rfWZoWaXDvogxJ
F1Eto2n87VsudRpKYdgScBnimiq333TCW1QlUDu7OKxUDlc2Avhxzv5WLvHcx7QT
DyY/a3AGIN7sfumbdnvUXzxU3CDTCYAqHuJ/iOfGH95AAi2vo0dhBS1IiQVK8kZF
F0lX3kqEtsIRzHBkx+BoR1GY/GxiCq+5OGpIM2kdUbtCxOsRjqAb9A+PqlR55QTN
pmuJ2tVr95APcZK9bCYQNgKx9weyRA5HIsrCsd5jx5KIPSsgj0SIFyTOCQ8sbfi7
Q4vFNynjHOUGBpFzzdM4yp7ffgVvxcZFTayg+otoFo2zfHfL25DI0Wx9lTKbl5+6
DSvjTZFISLM2DXZhAm9PwF38QlymdwEHEVkEBvfV1sGrQi42EJwAOKhK1uMON5BG
ChAjqpet/Pnf+CvnyndvWm8TrPIxrLsanw7LNdx/NxVmtUUQcSxVGHK9cpgcU6zD
GuLVIcLpe0NlXQvIWsEL47IP9kgkvRfJFh8Ybz6ji3WPkXmHRwJdBVlM1qXONQ75
5Kyj1K63u7eeW1xh7mTo0mWh1PSbvcNS3BqwFyNlPU8fZlHkm889W3qabIEcWqvC
WzGTcEBsy5Fg6dmtpa5XeSJLLk6dt9o91XsLZqSL3E6epu1SEPZmPC6ttr5Qqlti
NnzWsm4qqC3a4XKxAzRG4tcm8TZMFO1eu/16CTLH9cDuX/VQUhs4NhEnSDue2pBy
/6R+WUU112yiarxZUHspjX4WqbDG5CiakbCT/VmcJ0665H4APZfJmxPeeq0wOrut
q9o46LvWDtWseWNxpdMj0GsQcVyUyyyCU2n1rbBwswPgHWtkxNaylaEn7C2B7brm
n6WtPp9yQ6plG4FAW/OyrfMVtzKL+zCtw8GGXIwQWgYLdunqy+oJ85Gp31TKMhgZ
a72A/8/94TF5pdaRDM9/LkjCUCuIRULKmIEW5aHBv5B/VjUjlKL8CUcy/PGQIZJ9
F6buk8+jP0PMhDkhy1dieK2RGblxsghSUdKISwA8JJUPTgpmJSj7wS/YKfkXZqu8
r7oxXxecraBqYCdIn2ZVGVuUO2YotVuSMPRAF1Qrxjed7SYaDrIZesZ5Hd4kOiql
Jl5vVMIhD5QdsPdPSwL2uliD2JaKbrcv0nAk/49s4fjXSfi7xy+d10B0kmdNVqKq
y6lTwwWnI259ZsN5RIPq1dqF5NKbreF0QCoV3kFnD70Y1m7I7mLlHGctOpOz5vOj
a507FTVaRXPPwPfE5XNtKskQEvGwilXZsRgiYw/7giVE1DI8Vn7Tf0r77RxBaU3S
7eNBFub5jTdnZiZnb9LIlsslSmNx/nJ+BWWRXGD0XTWfUtWB9MLfJVH8iRF9PO5L
GotEN7yaBds7opqBApSelX5IXXRYc7WVjBY+hBGib9pn95vpo0l7gVoc11bOooQr
WARH2qaLrjDdHL89lmZ89kbF6k0cE3qKaYJnrTLdVY0pTqZ8/ZJOVQROfA7uLRJS
JTJcUmPk/mqHUK4S2cCyqc9UmZ9iQPFBC6OvliflwN+chIxPs/I9s5UWQQ5CsvXO
7/tkYVB6h5iOu4I4t8+dWfJRSGBEE+5RtiaXFXklYCkyXKuS2tUk96uMRCgR3riB
nz/y2LaCNiKDRHu8Eb3adBDVRLSB847hXSpIEsW+fmndD/YDPbLt+gnfJxCZWWWv
aEi9epYbNlamfcSiPtbOknEh75IFfxsmZCR6jXp8YmLXJVmea8+J9rd8YK28egrP
j8t6GRgpHclRRAbqyT8PbD5f1qljNbuKLTrOYRwKDEk/JN5YKvfMzItt642YQ5j2
l4WhJZmwUJHSWS53FFWmQ9Vl3EXwpBJysXqUjQzeplKIbhokIO09Vo+HwZ52xjCq
2a0eLeHlLPeD322tTViqO4ch2B/ZszJmeHUZUhYN1C9NfyFl0AA1MKrMjNKZTHII
IRnc+MDojqvLxQReffA5houxc5PYOQzfVoYwW2y2zStG243kel4K0XlT/x7tOL5a
GzXzG5/cKiofQHbQ9JL9PMJADGbHVjTtZ/wqt6Tfu7fIYqD7tTyV/2z7EY6GIyAe
p+btBFBYZ6vU0hED9b4EalYtySo9CS34mYjNAB0UVgRBMfVoSaye84QThKuxoqJd
iJe1T1QfHLee8q4Twmu6Clr+gzQTffoeBIsnze1PSBN4WBvVR5LtXlM07bBZ1CJD
6D6tEuNNpKT97DQFlDsfpQ3uI5abdF8bUz8oymzFJRBvmhz6dz+U3wkUNDs8OUG7
uQxLNswKfaagS65Kk3qUNRQYFz2JkjCeBf4+Nz0hAYmWx1V5/DfhwBPZL4S4Zlu9
tXApbfSzBxTnkBWM1kfiBy/6oo+lSS4pkacfF9/Na3MzB8+2T+m0kVjtQqhIrFwS
Jgc7g7QzCAmqiFb3MulCRa3tPGdLxaYVytZtIpuMdvCOf18tFnpqbfODwSj9CeRf
1U2+b43/pWy8Q+MNyUlEHYGIRGqE+DUeYADPspOrMYk7e8pRPcR4IXVD8Z6xHbDw
Xphg25fqxLlVYFsOxyp9n7yaK1rQX+Zk5HWrrdiFhBHI108NqqKEpkSdlhDpQjlc
dvSYnihzDm8dUd1Hj25q6c6GwZr1qt7QuXgjxN08uxVoRdV5h3jbClf3qt5Oh9gF
syC1JaL0wdPO7KoPqJdEVL2oL7nV08m0nW++UmJrZHuCkiTe966EUx8fILb16mEs
dMlUvysXQxcUV7gvw0xHbHxPtkVKEGvsRvhUwiSsG+0MLE5CyjkQw5IiHPNqpo5b
zegsj+2Z6sUMew/GPDnaPIQodUMQX5k8ZUDxWmeZva0kbv/yQykAd5FzMHyzg/KZ
AJd0BR9hb6C6OPu+PYibXWrq/hkvJq3ix/x0W/UmpkDBN49t/eCvj+zHBTSsjzbS
UfzbO8z3WdlRvKVpxrTS25vDFHyxEUR1gWyk0BS0+GVH17823kppujMWaBxE1HnQ
0c5eP+5ZMQL7h8qA8SqOm0+2fNcbDYAurA9jJh5HBRwB8fqpxvEP1Sc7JoTsO17h
rVJGKlilupxGGTKu7w2s3yvmHzGL0AXO4jvGZzsgt8M9jVTzYkuypIlaO0x3p30X
xS6ujL7cZlZx5PDlUKtcYQvvCn0Bw06achwAZak+dMR6y1lwrKxvK3zPPHHL408W
av+R7Ae/HpJpdeN0mRntic12iEVcF429AGgOYVHEm2uk8S3Snpi6U1mWnVO8JOBo
r/IpFTuYjj4ezqn3PNoDGhLQmmUZKhxgnbkYc04nYVdKzxY7uewLguGsSdw0YoPT
XuDUMttUCIEgyunZZ+/gQNn18hgBlZX3HuDhYZNMuqiNocpuF9fhPGxkHOu+UJFu
HU+LVKIuGDBep5ckWp5VIoiIWAyVFzqEj7Bs+ZUIpMqT2iKv+/x8M0yfjihKILV1
Gwmdd2rI9UADyD9T2olFWhiAxNmspFH8ygWnWVsOCp/5SYo3blUf3NTeIFpoxCUd
U2ep/On8T5PH7r2NokzOP/h75Hgw+xullik3wJsSR9zx8HtzGIyjO6ez8AQfEKMu
ldXw3sjCByEwTSIhzC8aWB4ChnfLYyFbWHwvgvJd1p8DM2PBTmOB+jkzlEb+RMWy
KyMoo0vSXoOu0KCfH62FVzq1P0VwSy+VwKZHiuMuHNHGnT3LYo/IOepW/1ZIGjAn
4s8Y3P+5cZQYSTzy4U8d7mkwAPPznfKLNgmcvW4C+/nFw8BEr5HwcD25qfGi3aY/
7wCQJGUlXnubNuK8VOOgTeNfIIF8hmx05WaDTZWM8Fea9wUjF5oOpmmNCljGRUSu
YNRP2w3/7Wq/20bqXv1RV1MYQ1kyHTQdCKKds18ATdRF8/rlmWYE1/g80XDQ4HC1
GgJgMY5F/gLLWSf7HaPdOUG2mskjFc4EXVHITOgAIexup+nKsC8736G/Vb0k09h/
mYpzt8ag2hE9YnYOLS/+JLWweexXkWK3UJw5pe/xjCN3cKSnIivBtCEn8oqWRGx0
nYyzdqO7r5VUFoS8JPKZnofFM0+p75MKY+Dz3Fu+SUI3rIuo+lftXEZEpU6B8wBb
gYLBdp10XY1DwuEcVcCm6WfGYJzMGB+xw04NdvLkPJt5400Eh086TTk969pRdD8P
Om+2qb54Z/ogpBHzKxzMuMNO9r0LoKHfGK+s9mQ0bKezjwptzbpHUsAHlALzpBMV
F0l6+FCbHSkLO81P8ZcIt1nEkMqJd0PyHahowbdT4vgOekPDKuyFwcS1TWyKuvnM
6SaoEEH4gIiTzfzsrZ4Ojcg7Flwhud64jb4mjgDWQj6/SRb5KW+/HZ0QRsJRQNrR
d0jYmJpa21S0kLJ2ui098T5379QHwOiR54FaGhaJel0/Qc4QKStO8H546cMNLRe1
WaWaP1Itnt/ndLHmBl+6lyxp2MmKK6541eXCSf7wr8FgMLIcoxk/0Nl5dViauUdk
W1o4zOYR8LFsU4K2OFWD/l5XELLH+KFVrOUpMpHFnmMkoDtE8uQKFm6Qo3wgnE7T
kVj9KGpWc9YlIuTi68Xb1x9DUusq9oIYmTCsTiEGuiqHMRpfXX1BOF7uJvZo4pgg
wjfRqG0cWZsavtnDWWOUtaP/gLPAQP66AY+21hlNRtKXnQ1TWdPoyNv8QrRLuQnp
atJ/30QnT5jPhDHckwfN4c/kWBffpDrhpp456dkNuV/fmWVShRKQKetWnjRjWGsr
aiy3fBWqeCikRKQF8Xzuan93QRWMe7WKzKR3LFO1wDAuMEzTyYfii+6SKd2DgVnw
nXmCTVaVwuEJNqVh8IDWaKmD2QisQ8FtJXY/9AeuEbz1ZK8PD/fEB9Q9+xpEp1yc
ksKhtooZgHIG+8CD2LLcFvUMDv7wOuiPlnilAghZmEBGXVPcHifsdSbzSV/l0I5G
yjFMzhrkDURw8E25KBhKXDkwptNwH9ejYCQSIqzR07wSbqrN7pZDz62ItKOh2azd
Ww76RPC4SwmLUdM+vdlaoP4ghyxcjJzwg5U5nCT0wvYLSfiz2OVcw0kmyTd+F17R
HuC+7osNuKBCbgH1hiAcqXuFZ2oM8AYa45F4IjVVtZlWDUPxECG2z1Bfv3IhMSym
vU+u7D3KhmMGWv8Yz1lkB2S2oFuxtgimjDTK5SAzvTOrnGzeWzhlQXO/cj0STic8
R/bEyTyuMv5w5UK+qRahnjrncztK1NNHnzRaMjja4O4Mr2Rov7KWDdyg3vMtNsvK
4k0ZX1xlRSD3WFzLJXpcDVVkmapEutpCteaMJqVs6LL7sHjW/UE1zvb3XDGGQBYS
zvBhy+KbjO1mlppFk3/7mQLiNsz1EaFQDju8TSvFlfU11dg2Gqvp4jOMdfvc5DaE
MVkzYSwToxows7hjrp5W9EyAXYRJW0AiOfdMCEO+6RUAekdmoOmKgcMy2j38YVoJ
U1ryWSmVIsbsBlf5IvzZXe4ZDwckCHH4jLh/fg9IdcToFzLahrMku/iRjefjjMD7
EuvqAZLPnxxekKjr23dLxOkO1JjW82DiSi1ZtahpLcn3g+0ymTiN7nWj+qj0yfjb
9+OCoxBWVaDyxW98l4R8p6Z7bCv1L9Wr+4BSlFK4ysMsRiWfI2DPiJ7uJvD4n8JK
ILtHnjCzZoI+GLXx2W22ca4vBTWouE3kaKAg5Becr0TSDu/k0DSBN33DvQ9906bm
uC09BMABHHxEBKEUKJOD+FqmwO9LmP9fOPmStOXK3+AfHGtezSdfK6NqTricYVKV
W5+ph+Ohh/IV+9Ap2KfSYuMGSxcctZuxEsGCs8eRFmsF5jyF4RDG/5PxE8BTG4K2
WC8wIuDE1/qykf2Fe0OYIKz1Egeq0AZf+c7gL5bN3MEEOtBq2QLtRX1b5ExepRIh
VS7Fidmyi4BH3DxHgrdK2VEpAWcdaOHvCR7HrfMV3aWnZIlGlBcd++aGto33+Le4
kdHX6Gf+80QE8WWwvCOhgYYvJKbO9kiC80cfP6Vfa8Kvrx+H40+VxmJXgbys+YJU
ALnOLURXcnNjEfW3NwHEIu5RsC3hyDhEnG9YQlbvhk27LjxEDsbsHKGJlbVWv8wk
dcReGtEjWHMq52dzlDHSMjQzGIkeFUYpTo77+tJ+doqLSQbKvg2GDsHH8dULCIZB
cXBCHH03h+7vu3WZNJOaufIzWyxoEl0djGYpEuekwFsoZDtixtrlKF3AP+Tk8Ino
NnNEbscGvqmjCPF4O41x2R0u21381appZ/SC/QuoWMCmhg6M0BQRKytw5jYMxqtK
cadKUCWVr6EedZxeqin4M2Z/Zo7Hb0IcGap4lezkxtZkDuVHUkFDfsYOr8Sj/gS+
tO3wHI1z7DS0GHGnfMOSnPhkOsoNx/UWfwez4Qjysbmktyr4trj7UVzpfFf2oPQZ
uHRFnMChQEODroarIycKLaf0vK7mBdUAXR6BbDMB214Nw61qJF1jbxGdlDKCalea
dES4ovwvs08MgWkOekkjh4l2857tihLGdTHEg6p0xmlGqIwB3onKtu8ADPloKRHy
KS5lKNwCUA6PLnDZXvPdK36kTwj9UIFoj8rd+AS6mYGkko0x2viBBSqmEaicg1s7
N1a7vQ8tpTR6s7g+KhTwhnqurLpDTkt2cI6fdgxMXsoBx3DoBThB42Skdc8G+M63
4LABZtkviP+900ZQR9wK/qKxEKXTzc1dQOc0CHP2Ap8qWBbIPju/zHQlvVIyLfc/
dT7MFscbvCWk8czm4YOOXo6FxQw11ttn4nd+qMqzz6AdqBKPyOfTcg/50Qm21Quo
bkmWcJKw/nxFqA8o2Zw60wunUDfk6Mxx1nj+Kc8Kx0Wm6oqcbfTasocGDcbOWwvh
nif5rLRoGq0CpivRkLFRhBUJBc4474KrKHgEsHdx5TRv292eLU0Rcnt6Bkxu7Jk8
l+dadHtdFuOY5EA3vz0JLQaCxabnFVOpVrWNJgRdRpyfODitBQ4is9l0p4eg8vXN
cRMz8PY9QDxl+R3ztNOYJR0hj/QuJtTM0p9qgCJhAI36m86nuTmRLXUDKpoJAnrN
ACfTj4HJAeFzou5EreA17td1t5Zl0FnmRqz+hD0Hl6Lo7khxv1shW0bz/GrJF3Qq
DfkgqkKaEy+zi/zCAbYooaSpZt0sqz8DWDNE9f33+LGUtp5GBv67S4O3UoQTcjNN
ckZCfT+7QQq+8Mk4K4SLoSI8L5x7skhc/GsoBKx+QmH+dJnVAB25mSP2NbVG+sLS
PZmUb2sldtXsQVCq4wVpLdrLTPzE9pt7VU6ssriof+IydxX8DjwxC8d40DjIO1Cj
sFbdBYjuubNkaLBQ0cW/UtKqPTcwWfpagRVW8ma8MBIWa5QLfFlPndLtUjYbLVmn
g7ERsVKDmpEgwDwJ4i/qMzXy38T3yBbcDAq2SlUh2tJqgIftJq1X/HkxdGGxw/FM
sjoVlLdGcBktJFXBAWO2jjHNwZf/mqq3kc0a6S8esCvpbc9PBr5MONGyWZ+Ye4oT
2v+1VRSUK3/56Oq4OoVYsftxh91zBHF4Y/D3KNT3UoA5qf94C8oEZJ7itjnmewOo
n+v0i6UGijqLAOgW43AKpAUxqKeZpZuOedq2iCMrzRqW20gfa6tsp0ED9mW52tDj
Yi/G3vj9o3Ey2q7zIFjBVlcpobR3wWmTQc6ZtBhotHQjesEHMGImmZJ8tVSgGLtJ
rJNtD9+C2LxqZPQoyvw9rurUCtGxxKbT7ChK00dxxSU52LIWWfO8xIcc5qFgJzaf
2D+8FTL7QlDnzwi1n3DtXudjB9MGXehYtly6/xYa6w02Ak8/IrqAfLaQbsWg8X/K
yZ9VaO4HMDm+cjpt54ixZvt+SGEOSyTdG0erv92gl5hwRYSW8sUzVDAq8FqD9lUS
KnMwWowjCrA8OkpGXniMM4L8t1bsKmnRdW/kEwwXQokVd3KWz8cAu15CHnCTuDbQ
ZvoKoogsMI8flH0t6hKJjaRvCuzLSr0xEzz4MOiQCdjTYKS+8o22xhC6mX+ytrag
RKcU4BWJT5AWKHYHc5VdQqyKGDonMotbXiU5gKy/oZNNxOK8/XZgPH36HTGxs6Ai
eHl4f7Yc662LbrbXntcqFc78uRC7sahq1OhD1NxNmSWy1LWO3iLQlDr6o8qYGxei
9AZb1SxlaB4psnpfYt1EBDTSJUGx5tHWmdgLJaO/wrqEi8IFtelse13EW+n9tC4A
fuvgQqPTEf0Owg5ao6wD/8/sQvoMOsSfWYvH8Ghpfvwzqlqcqzg2yo7w5lg16BeC
X3hVoe2yoRmm39N8fUQgwyGPn76CYkuslyfblUdQuOmYGKBoD1Y5zUVW1cn7M/HJ
KQvCBqPZJCzv3eRzOSi+/SlZpGuB+I+Z/zJ1P3ZuyUg1fDCnuAO3jgZoXX/HqFtu
eZxnpBa9Uv0RN8iVzBKVJtDmDyh8ZDB4zDCtE2ilZfKDkZqqR+p78KhMNBI8bif6
FMdXvEcQ1R3+EIHeTq2s2axiFlnwUvT3W0e9U/qPN8YinZgH9STOYYKzx0FKMRWB
r0mXukc9unWTmWrPR3gFQPGdXdj0lr9s7iB6ZA2i4YJXJdyZ1ERpFPadLnZdROZ+
je5N1TjxskFgk/TvDd617mwPfJLpiMsC0dVIzUB+mVA0F6IFOAEM9XeD1TPd3SN9
HBGEreaz8iFxmX5dcDFU1HfaXBS/tWw/P5t7RdTPAYfyFb1Lt1iAIQzKRjyltJM7
xOzhcilC+KSl6aW+ktRprSdufb0Am7jiWVOHON1/6N8YTtxZn9sGPb1i0lGAl3s9
RgV27N+F7hmHN5aIUywqs/un/IP7KgQ0Xullz/bEdJJ9Leyu6zvv3mPhWx+kpgU9
2cSLVQSvH9DwsyuiXK323Cf17+INuiNLNOJ7JSOOjLwzNgnBOApWB0iRIiNCojwu
mP62DO2XVOjLc9yUZCj72VA/KPKgi/OtzJpplfDbKHkVK60hbCHIwB/j3I8AdhBZ
FnM1MwtRpfII5XJ8xY+ScRTcrptbewhrq3hTRveaEnxR209TxIQgzi8kQgAm5YJP
WH04ujVWzwOIbLM99Py+ie9KkMvwu+kYgA80vEltHDDf5NurHi9YiJ1uJNwMxxc3
1fQ0ewu7oFM9DiehthIRRXqOmzpErta8XSVUj3ivL/X30wPHgzBtbTcphPggbHUZ
3Ev4I9Dkr4USyCOvJODJ84qUN+1lIayNH7b/8A8FIbyjJFLJdou15WhKrPxkS4jP
rJslt687VAHn0HEB1i5zFIBLJQ6M1aVUcckj43c5dlpDfUm6SI0XFAg4odIVGPls
hiCLiFqLhLYdyeN70iajJwnXks2c3ODqEtDN+3h4wMLoZhtmaAqSS2Sscq5MHa2U
FJ6kZc959l8JcxwCU1ZVcJrQPGdhb8TBJt+BrtN4ziA/9BPjYXYhjx4siugvAKum
87xTLdrK35cCKQIsmZIhhkx+SG3lUZWjeAziFEXEdOAJ2sH/QKa0S1amGpKgL7pp
fMc3DNOthnR7jT6V2GTtFTn+62iDQ/JyGV6rpNarjF2Ouv927wwZOENrXa1EVuVi
lzXjGQ5h7+CoHLywaDKeiJk8Artlj7+qIyqshqAJ0SZ4OLoOxDpEBbXrbFwHvtZ0
3+UBziLA3wxRpDduHnKhzMDjara3tCPf9DI/cSRlnciJ3EDketI/JIHC1YQq+bC4
zJxkW+8pW9fxzwAzM2G6Np8fDU5Kce80j6qf985SGUXskn+KfyuHd/lGnmxYsQTA
WyoxhNRSbw2nKKvFwEBvsHFo/Eh4ZPWrzyCMeX2PwGccT8KZWGhSCXW8H0cuKn8s
Fifs3U4xtTdykzvHRpuYRWIiVJL4qsETdlZKTSK/1uZKJMY7JcE1BJShpcNxBVP3
Leu7n53ox3h45zYLhOgOq9x1zviTd2FmB0DfMliGZZA6cpF247e6WoA7tC6vS4GM
OdsjcXEhGu9fffO9v+ngVC+TF7WeyPwv9j+YwJLL6CHO5bpymduXb16VY+j/Wrx4
y77nyTOTxIakQS0b3V8jlF108+Th/fPWzITBCwFHZb66XWMa5n5dlBWE8d4Sgg6+
e7nlAXDs0Hywup7NpxTOfAGZWpLNRzovpCPbfv2ekUMFSPJ/wdProKV1iwIhMyQa
cgLC9NLJbDhEBSb7Fiqc8Go3nI2IXM+95H9YAd4X05hQhvUwoD8ehWvIbQJWYSFm
e56ndNNecwz4hlb3KiCAiUPfLyWFP3nuhOUE4NfKFyKj/d/xohYPeDNp0/Y4AtgP
IOKHTHjag/tRkuE4sKd2sZgyLT8dpJ+BajC9ABl7igmTI7FTWyg6Rv7K/Pd5vluL
uijbOxv0Wo655sYGo+7ZfGLHraMZ8YhOY84NObJi3H0xjM1+aCbJ/ncNy0NrnkY4
BvOk4ViDxXhgOfFuVzLf2TBav0tWwbHFPXzgWo014oE4Pcx5enQivKDftiEhAZk7
4nSilDydbYi4AeAZ4LEC5HHYVo39Mx6+Ysrb0Au0Gr5fDQatersjFU0D/b6phsdb
F3gAhDroM8wMxhTktFuN3H6l+7vn9MCRQiyZw63MX9/Obmy+9ePOr/hXVgKkded4
kxZ2JDA0Kdez2GayFbhjwXigiQ+TrmnvAMMxEYLHrD8hvMOrPrCdBCC/0ECx+Q04
s7vfoxttyehvxsH0XmnxxfQh7A6wU1Z6TX62ZTtmBaL5FEfGtIFN7q3y1csvO11H
FcKL8Hpl4wsi92uvDb/2bKgQRD4WnuZcnnbr/XQa5Sx8mw/6JDNQ04QbVLuLDsI9
ddBDFqj9TQIkRTElrCS6D4EAeuSFpzTGBmrFgihJXyZdKlqLiIZQiJXKsmRU+SwQ
1GT809b4d7C2pEMaduWeGl1EU0m0v68n0wKL41KUUGZuykU1cYcXtHEv41Rz0YY0
LqSF2c0qoRzWR6cPtkyUL5NERBdUxNj++bBc9jFKGBgVjNrKcILqKGKjcw0F+TGt
hJJZJDcfn13dTvMMJeAJ+yDAPDRzN8vdUjpiFwmXcU25Q85SeKDB3SjHW1D+rgy6
cvDpSYV9yhM4XjPmRZTI/1I1DScmIY1OQFZ9GGb2hPkRpNK5ta6NWbz1tLPqZBvH
jGfzl8160qhYXUy4/7ssUp6b5EKba1L9f67uZsUOW0EnvmGN9YsK3xBY91L7mFTQ
9iz3IsjeLBK6RIH1Qsaetw3JxEkPVjuYFzmdz7CynZm5S+HuKvqKeEAXSdF7wOjD
+bpC0hVf/2fvLGjwUj4eZ+PW3dPTiuK6yuQn7vj25sTrF0zm1UE+x3r8L20Ay/Xi
aaVZ/djKIIoQOXvmGxqojdfC7GDPYDCMPqbdoMY40PYdW5idGnMBrPupK31LIebm
RZgTgmv3wWV99OtAwZslAVdel1RAGF3mdeK+JP6hOGpuVzfLaY7ZNk2mQackprne
rmq06C8tEzMD9Tg0Mm+nQIEsgFDRnDFXSZQQUERlUTzk6r6EAVWKto5vE9CkS0ok
yCf0/xvifFUozdeILWqAzWhub2k+3u/7qpjZJcERFKEx7aJKsZwh+mnKawHLX2f1
tuWhDYYpPxUQIE1cBpZqDHuX3Rz3LB9OJYuh0aR5Xi5bocwzZFv+zANiQLVxMFSd
uJwdy3KWLLF+8MKW2Sefi4EZNZMgHMHeQfJrzEzKbIXzeP3V2Srel19unC8j+Ohl
IanwoNyRVWuoTmGhtVjHX4MOvyvOLomiFje6xoFb9JiPoLKeWT/KOfoJJOqGyC5h
mO/Lw5sT347m9iY1lryqOq3Z1eIFZoge5yUXP2ym1Yf6hOlPEvf8qWqeMXDg1NZB
i6kQtbBkI4MdZRnaGCBs9RcUC5vIZQUZK8L6nY+uwBnJyFhrkvoYQcCPv/X6oScu
zQgmkadd3lXG3Lpwduvy3s41cVjr8HgegP6QQxrpDlmBjQRC+yvBUwyUrpQi8pMj
oFEQ31fFdBXX/YS+IfJHEbIVgaXZ8lvUfRBIUgKJzSu0ANOQ2OUkR3HhVUTIL9Mt
sXZvAWClr32yV63h3gLNUgR/P5yP9AEINCHR0S7d37Gaj88/6aCeLXp+n8WkQJZN
c6hlDvx7Gm4GC94Nlp1sgK5YKjYRtQp1K2sQ4uGLhor8/MdSwI3/neMEOtI7JEQI
1LXnyzmyBJPLCAOvkuFTqBKoX50TBVVdXv/wgx0ND6n0TRWa3eHdd/wbBCBC6cbC
q/DyxdElQ2AKK/g3v3whqn73uAPcsrzunOK2ouGS7S9jD15p1MDlE+u/SiCQtTNo
9dxRxTLmeqWjxinwo7AW2H1cNYIeoeLQdftNBYQtMqPcZDFcdqgOrn0xN/sGbOnC
JrQftPWB9dIx7Ob7SWOVCKdsVU7CStpvjNUtisJpcD2/40QNpOghIqzfBaqIuoqB
U8MAqrO6H8lm0NPwYcdMmBYoXNIhBo1IZMIZTUOkwHFMp/KKPxN7ORy/hGCOVeNp
fho9DuXM+nKZTNkDma5Ux1JKgCAqRr1ejcdVmQz+FTRxLDjyKBXOBXgu4it8fPCR
JJ7V59vXuz36K1u0d+cPSw28u3KGqBb9RnAEhKnEgoYZEw9bX9dEv/T8c9l9s9r9
B9GwuefILYFYm6oMwUBZ6kOrxDNLCKdO/w2bvyeHxX7KcJx+8NuxZcOWUxwktbaL
E4ayi1HsnDclvFioQarWXkXXGlGjy27vNyS7xpaSeSByd00Go+cg+FdhYn00pBvG
8ISVEGJf30qnqvFQJtiNVcELyrg9VAY+FJqj+oy2TnOVDFaRQwKo7mI1qXEDzdRv
wL9RTq3lN09xGr6q5WxTZSrPnZNpFkKtWkcVxLAU2gda+T5qCU8aUNBjGLsWVyvY
NfwGc2svOhINMyBEjLsT9R+0t0wl6XHn8Juu7t5IUlhT5HDViyJ8zUn+P3qZAGop
WkgM0d21V1ndz/mLXDOTnsNWzMBX61sCTUfuOgNLLiYMwqVAmm5rWh8rXVukEdjb
HJlpCR1tH4FrqwDunZvyNmnbdjgj6OCeACUwpXps8oIf26py4bvcODVA8fI7OTR1
bBHSebRv9BVeZpwFgQS0/Rx2helJD7CxAH/Py7ytv9+FX0rm9+1GLgToc+4SbwYD
Jj4pQbHT0/MXQKI6MQ9az+dtdkMsjTGm/xau/joNasAXFcWIUk0/EbJtiNKYmfOg
AEFu2vKYL+dZanTRAwOFtocgAEW5WIl5DngJvpPyJg9tDYl4r1A3cnzqeIA1LqJD
X9Yij/6ICUl8Qv2YeeP3o1F8kPcVcYgcPIxd5ffvQkTeQNbzpzwQGqGiXDBuqsck
cHGsh3S66HNr1UpH1xuvbHpts8P5yQa3qQWOmM4mKCjOVh/VyXF1oiVn8GoEF27K
bv1j6t7++y6hRR+31xYp3kY3BkD3roo0XitkFV359GvEURb2iZv/5Ah5Sp0aGi5V
PEQuCx8cUFI0GF8tiRl53rJAngE8zicWter2v1yqFdd4FBTtyJzDcCWGI/CBeCNq
nTiP33MhGsV6SmHM/Tpk0E8fI7MBNcQgMFm9g92GKb4dlM46KtxbYvpMj7asH/pJ
lJdo+CvXtMJc+hQMFSk5PKbNp2+72uZNvLxfk+R1Eonyf5pOOxbI5hEWB3P/0vWT
k0BXkNMULOB1eIdqvnNpoz+SPvx+SCZAspZA5Pcpf58M43PPdhhoVcD7dhAUXE2c
pLCou/xR/7gHIk8T7Nte9HFulkPYS5ARR5EQsglWcv56a2bfGXMoOdhSbq1T00pU
6WtHcQuwZw+bM2jrb6NuiGIiSQzrj+XYfIKiwMX/atZGjoBBewL13jQpyU7ptgQw
/1KCQOoslWCm76RIDk2MF7CIBE09vFEdGvYaLPZTmENIwSumV+BjTjfrlRXNhvTV
ft2kf1YMG+WbkNJk2kj+IuwBEsTaA8x+ItkyrPgiYKVQIC1P/MQRJpC15yd1z8ZL
T0ZtdOffg8MEjj30dzd1ED5AxoODuwZF1NlkvdwPxTBl6kIDlSlqeDCsLBGk4gjB
YR44A2xHiBnWi5zZgUww5WMJS5iGuqwoJHvVQ9sBaoUGhB0vie+2JNMPz/9MkPxN
DsPltf7kOYRrhbeZtvMCaCaXNulobGhCDaUSrexCP5j6MumCoS0tXz8iIyaSFITH
3QaIET9IkB8ygtO01+XtHNXX2mwknkkZfwzobFUeqR94BFtpdqLT9JQ2gHPDElxx
qWuT8KsWKdez7skr53qQyG/gZxzBuf9Y9qVuPVzqLBQeykPVvVO1h94ZALYUyo8b
m2zfXearUlkfOiHCNQ13jrd5Xhzcejl+J4Av4psd6ro4j2ggoeE1X2z6VSTjmZLx
Z7scp7B4nOAGBjkgvyiio+ijGFZV9GTt3YBCkhIOuvPuL4sxrFmXoCJXGK+hpTBQ
/+pn6fY37BUgsJmVKIJFJ93l0zoTWxZTXNJw/KHgKewQvjBikQJ1BLKsHmAl7m0G
oq2Z9WOYkyzPmNiTthYg+u6SeRo7y6hS7APir+Fez++19s1qpjrfujaAU0KaGEEK
cjcuEH0Y6b1lRwlhObcV3bmotODstTAntbpSyIamIPIUeHog6xr7TKtM7DWr8LE3
C7H3qQPlY10xdVGvgJn4H22CVO1GWOkE9TbGpNJytPf6ukWlH5fxOhnDlXxxB6hs
qp88SX+FKAYqfYg4hzoc9EnWCPXCN8T0v3bQdXaiXuOgEc6Ja6I3JGLRRIYuGjid
Af3jTn0Kz2pTZjl8LYUVqm+3KYxBVTm8er7kgbEUhr6YNksaM9TCWbhWWMEMZsty
Ofapmb9xcw6gbmM1IK2KMzVrZ4DHcWKdZZGa+oXIustbDLCN5gW441uh5aPL1W9l
hLs7lY6BHPCbug5veJvfBh0LYR6lKuaxsw9khtutyh5Bc8To0FgjgonA82wgYdef
z5wV+YLuC6ovemaqImV3I9pndY/A8+TWhRRoonwvB+5+uDo/UFP/3aSDePuPyu9c
rOQ4F2UdI/HXEshwhJ2AGkNW6/n9EBSrDItrrktn8h+OnotdR1U5jgfjhdWVon+S
tA9glZzLcVSDRNegsaxJBjZosZv4pbiZ6s+JgaJmfsAgr2aXPv2eT1IipCx6/vRz
rVWrE7DBYoF2TL0+C8EvbVq9icJajrlUh3QOU4GJDy7hPAdPUpM7j3Sib5AHMR7H
ZFxcO2k6Lbn/ChU0P8y+o1fqfZLe/gUScHngBKQ7gZqBKIey3FnrjDjrAe1+/4Im
8eMwZbdZxLjVTuCeGgHt0RbW2TpSTyCGYY7CFXVsUB+cAMPS61TPektIhFtMBQz9
uzjwvp4omu1RytDWUWMWO55E/c8Cq6QgsVcMhriHlLv7N5v+oPXTTpQCszFG+PW5
cNcbKtj+FIxr8S+aYdziFdx6wwEA/Gku3Vdufv618hNXniRsT+MKgTw1hJA+gIbU
VUrdma8pwPVHubzV35muzBaVcUu8OPRloogq5GQF8hVdIVNslO1XUZGQ302kit/l
B39/BNWuaewm+JG98AMF2imho6WiLRZrl3BgapfKyhv+bdjirmLJVcFW8wIEapC6
KTB37Ak6Ey47wBMGNXxI3b90Z2jd+sw080uQ+4T2fZuFyTc8dpEsQ0XzJjEstD3r
6c7HRxxAKxur0fWC9b52gY1TS4QEKUp70d+Ke0IbbSGck1ccSJspusPvUirL8N06
voY4/CzQWNhSd7Y6m8Rb2MbkzmWKYcZ1l7UNEM2WWrFJtsf2+MoImhfgBjjSch3t
CH3aKR1mJTDRDZ69A2S3X98JMx/p9fvUo2NUmXpSn175toLUg5qNrRS0USCyobLQ
08iCCKj+h9PXjFGlBr/iIBaLga1rOc/iTkPR7P/G3DBznJN9n36zBkahyuc04Svj
PaNvCecb4BU+SQeWHKMY9/HfWLHRL+r9WuwNZQnSSuvpkH+fEMLLFJml2O4wxV9X
3UvKOvyqSf92A7QAQ0y9W0a0sJZ8eHD5E6ok8zDypO783Nmt6XeNWJ8W2cMUaBGp
+EP9m3eF5m18gniERXlqxSkHk4O1ItR0IQmOIao/uD0gYX//o1NWLpSVpfZg1EDH
LPnpU9QFsmHa8PJnhz7tpnisKaVFaNHdP15ddd4oG1YCO5vsoawAmiRVR77SozUj
mFVSzdC7KgYyO/q4mIYVb7GCsYPnRQ4jj8dzFn9bH28xUGznkUQq54KjwGNHeGJ6
GIMgY+dNW1T/06KEBY3HVDvlcCo3zd2zEFcrR975Y+GzRu9GR7eeixyUnQErtqiG
qJxc3C/j4lj4f69l+Yd/7He9gDQIUvxpPn9JyaRIp6saN9SwaISUvpGz9vC/JfOn
1J4eojoFAv4FyaNcgsvCpM1QbVxIADd7Q3QfKlUdMuZ8t0333Gg1L9T+r7QGALZE
FcPQc5BI5ohEy0akgafmRCdWdoxGb1mRkx59WLnlw5Esmk+eK4nJeV9Ltxlx2wXU
DU/hs3sgMnzex376tqY72+yTN2rULVqml7AYJ6SEPASOf5L7USmzb3bI4TwLQxJw
ncQNyMNl3wg1zlurAncFd18nNfJqwAqpEcd7Ynzv9RzFH4DrZlwv1ZLXplynWqNZ
+Z7+LBkYGXdzpwSIk6l4jjWzottFCCdWu0GSQJKGOr0NTlDZ6oV6K/3o71tQOxpS
A5/P32AHYjGPOHDP6ftvMIkcm786SRGtAAZwiza3kcGMVzYcBB44U+ZLwe4Y6hLk
qAAa1dfhOxzsjS8PD3l/eNIxZnqY4lekngsRu2rUiUaBAPTyL2YW6HgRQI3wyD9L
2YE8/w4LC1spCO6OvP7qVxzuTUDn/W9ME5Zn7wd6H81PoC+6j/b+u3P984t68yTb
YdHDnLDlMb89pu0usuoSxfwNxB5eByJscnHL8LB89PqMKSKVq5M4aRyZFVE5ekOe
a0wD9pTPicZlz1ue+r6fylFEGzIlGUn7d6EV9lKeTde7a0ZPIULoO6axvNQSVAs2
OlSta5F9/0uESYM7FojdsMKhg9D2gLzGWfKirIG1R9V1w+8Ao7y6pV0IyuvAo1Ce
fG1I0c79/IcLVV3qQMsv6hrsqdTCEzqQ4E4kCJb5ryiSKuMLjiOWyLF0ZVIAS8YQ
gmgJSEVVbvL/zm7QckcD2VfR39xlfze6WmgVy8aM1p3OHaHazNYIJKQLkfBeKedv
tpQCZEILP7IYfvfxfzpLomf6wEhTSKSvnFTGBiDUUxmChHmIk3n+9cwKMqtT0sFO
aez1Y1BAQWoOevZOzSu7AHtgpwUsWX34lwBgbC7TjducQYE246wG+tu82MOmKMFB
uo+uEevBodNeQwiKFdh55uGbpp7uxwHEJode8FaQMCniCER8o5X1wRGl2fzU/2U6
5/BTaDqiXu0RBjBU3XTSEgpfLdTi7YR39S6+mNUMWMMNMEgyyZZfTbC5BfyE2rqT
HbAvKc7jc8E+qvi9oXeuaFw9YhfI+pxMzXFHr/3t9QHaflhTOrgXcjTEEBu944XS
g0GVbhZkarYWJtX2C567DljhodPyQa/UVQfRdwzHpC/bfQCTpTKGv7wmi23Ug4Ig
vtXl32GoqrJK1q/4pQ6Pl4RUQixELgRCzzoTl1rI4iQCdO+ESIC0t8gVYOiuS+J5
/BLGDaW0JgidlifzUIPO1F7OIfEpSj8RtmINK8GUY3FPwEWvuR+nMEeNqxEBRee8
6RoXHuiAMi3eE6gAE0ivtNXZN00avqLbO6WjGHHY/fBvIc0Ie4k9b96ysYBBGVcr
ZYs08DSg7EOxVdkWFpFfpOCp62ZUR7XI7Y4Rl5ijkdYR2E/RPGjn0egPj1dTuO6+
YIgeE6npzjUjtqbTQ9Afco28X+tss/pwjpohkM0xCDMr3UJpDjDv3uMxQA/Yyjo3
TzvrF4PMSFQ/Fkn7GjSQRx9Z6KUeD4sqB7qlns/RsURabEpTZTWQd4vvp30lhSNe
m3F4Sjned9NFWmTZ7I+lEcRc5JkR56Bdy8jqxaqEhx2J+r5y3JdhO4PS8Ps6N9Th
K+uk705zT2Aq7aW3xh+IvL2g6rrGhdfW3geKmbDGibXIrpCLWhi+nBV+0MV+ZrFQ
Z5q5cdHkIk7ZOjhw2hn/7kY2hhuA4uRRpcPhDl2y96wwwBXoyYW8GGd6i+VPvpZ1
qxBsUBedLgeuXJfOluokWfPjrJQUlGxPZsXDNecyhnXn74F4Juj+YwIr7wBF2ip9
WSmqMfnVhe02mCzVlOqpIwC33kOv6WijWjcOkyhgGWUTw2vJa/yDhHmOjorFI+cd
uNLDQ3H7bHygYTEkE6HiNPW8Lqhwuiov5nK06VaGyGb59H7QmpcZq0qDt6lB/J1L
LwQ5duWT2jDhTnXjY+UcEQgwaEpIQO2U1eLQc6b1gy5vsEUQOybW66KGP8dp8Wig
FO8tA2ZSvwGzS1L3a4tRazwgzBwS6KPVskUKD0RPl7k6zjxKxYQfTLtn18/VM27l
Q8AMKj8vN8sKmkJsY8Z7lxkRYrpYN9MGor7w4k0+N1Jgj7DkYEsBNA5xXNsFa0cA
0+wXktf+vLmvhf6ddDhJhfI6sDPqn6rxIy/8eqaO+Y9A/F+hSrWTMz4OezIpa74N
0LSr4H9YkwDBWG7y4E5ke13CPDvDuD/eC+rpCiWfi7hRQZiae5BT8Vg/loStVM5E
gzCmFt49AFbtjWeayMv6aW266MoBOM2UMQZtfQwSLAiSLrJTP0/k8f+g3mQTvGyw
RMgF9HtZAmlE/i1mzBnkbjJsPF/hWQlJdncC5z9U37ReEk8L2Na8iT2I2kfJDQaF
MxI7cXGH4In2Ar+LzekzkyYtUMSmmAeGHGT2UcXyutHBktdaT9/fcT2q4qQa9YEi
CoGO6lmhbQt4CBK2S6w1+RGudMtENBv8pyLK74BYCVijrjv63hwmVzlTFWHOrHuI
hE6qcEgc+ZBVhr+QdaOMPj3tzqvINAk3mrYjGP31lvjZ3X55qldMNSIXa1Ux5de0
UXcdChypGk82Ck64XsWEtgBEucNu+hT4jLeAGjNnKXbH25EWbYER8W/imLBGkihY
8jkt/yTzhM4es3eWtaUSkOf5o9ldgRQTO809qcIrhD9i9Cz3kwlycm70vcmCeorO
Zf5ypSsanV9jWmTPuFyMIk61IaIdSr8hQbOW1p2Pga6/ZiFRce+ryvZNPuCFe7gM
a1BvJPVe9wYrnSeyqqYSynWPK/WOdFthZNvN+Itk9AhcTTYdH8DluOHZtS8dzChx
Z2VhCI532zF0VG5sb2EuTWOBR3q37dChXc+W7uEMwRSIyYemLX3yHCnE1VUY5Ng3
mLDsvGHY8XGyCmLzTBl57xPlM+eOTcy/G9P5oLygisEz9BsaYOM/fi52EyjJNCML
phMXDqun7m9lboa0JGMXeSR8zvwfyvYkmjTIcZuYBm6xgfvlXQnUhi+4ZVcN1UnF
cjlKJAeTOab9Z1W+o00rKdocOGI6gMiXBK1jLGpZteIN+1rN3I3k5JD9BQDQwWYF
k0VwghxrXinytfyqFF+0bpKsySUuQiCj1xlaIOyTFmhgz1VAWejkqsgx0sxU+MQw
R9x/evS7A5hH3zCyVFFJ+I+e9H9ZoGDPRArXaciGzqVNwcAdUOIaSF6XJxlv21Sr
4E9wGx0ux533hv9u+w+C7dSE9ytPuLwiYyvM1Zm4eN9A1EGdZZNPtEzpRdEVWMvF
UHCEItNyP1UkTzCbJaCCgyK7T9S8637FFbTFd8bFEjS+XCtWr+GUlLzRrElREiTZ
IZ6NcKjcmo9VPWXo3eCvRSEfWxk0kTxD79DBvxV8mLOz0Gdr8dP444rkg4aKjQhX
KuIDFYH6yfmoSeWuQ7SbH4NMahWBFRjXVa9l9HMbqY1bas1LFXEOEtU7AG4DiFE6
jHriYLdW8EG531nEHg0FLSUfoEiUMgRKz1N+cceh13ENw9pFZYrCt5xbrZ/gnZdk
bsEXHMyApkVStF1n2a3g/wiv3nTiBceqaF+UqrkKUv8Cy2NMwh9D6G8E/FQ9ijYM
+SB2xlDIR9AGzyGCrQ4Fey3pMpAN/jOXvo49O8d0lXw/cAKWtEXNj30l+ECmSsm+
phHux6mYUQ45LJR7pKj2mFX5x3P5HHWbgDwsXaDoCd2vd5+d2Ipkarvw9DjEjMT5
09Wp0xQVYcY35X3J0o+iiZP5NKuAr4/DmQjdEdl0f/klA7C4v/9KNX9jFT5Qszca
7fM/TBU8umoZzC2MZ9HIR0IDy0n3gTwFCShYVqRhIv7aS44Nyf+2kDOsVg4y5PIe
z3Z1GbXzbBYTAtO2cPVYouoMsLW0rQzE1Mxw1mTGvtO/uNpoyhkM/ce2s0Akgx6U
PzbJTvfZx9iK5lJU0NJhMQENnqExfQxYCWWInoIp4khqIRgubrUIBaFs6yj6/WHV
zyjfq25S5mihpGIks7l3epBTBvAmAxTmomH6lYM2xu2jjnFM0kTRbp3YmM+PQm2E
DPqQ8ztF10+FYvySsC43rY40J6BvK+wzGUR6hMFLqMTifdp83jqHkOOenhnC8WuX
zqbh5AYwqcnwFfZhHB8yR6Lgke1roMRtnjgtd6CS7YE7aW5LL8TfV6Y2hK5MR2XZ
zAxvZzhCzVsD4YXvZU/Bn9izNJHTxNnuLaDJc0y1yBiWIlgwbrOrUIb96g56Ve4p
ajb7XRAOlGN6AFGgJblXZqQC9QAV+gpezL+O61qAbqoRcK8UchBLfRsShTYW/IdX
v8kLapD/iAFz1amx7oOz4GwKDFMtmDWNKcqOIADRpGNwCC2ea4vQ1s6K+52Dk408
CDGicDsMUiIgXXNEWKxFjCVR2H4j9Nh/mKg++bNBnYf6K77yvHMyy0qDdUsT/gkt
AMXJ3X+DUvI0bCpPmM2VDyn2afLjKbUWNxoWs09XTN+ex/fXoyC8/bTCX0xXO0v4
YVNfUgI8FPWZD0rycetMMoyCSZdKijC0uweiTxRyx90nxMb18I3lbi9Apb33/YGj
erTPomOoZ40+PGmCkZPtcvsXvq5W0mDDDWn/+6v6WJ3fCovQ7tQsyB19LzdCZOzW
VL+2LzA6R5aOoiR07Hkoqp1Q1w6JSnB17IANFtoNmm48s1eq/qGL0fRvX32Avmtj
odhyJ76sdGQq3vQvMSEizeiYFn2iunAZ8zRTtFZTVkImDvHBg6uPhgws5j8iVSRP
q/uLTsfY/4YGY52WxJho7LfnkUHR5T183++YwLxXHWK708NVfqzCBQ/grmfjYmbt
WRovJFNW+pZt4Mi5vo3PGWRC8hLAvh6f4TUPsrsBXNA9t0WvBzuqw1DcxThIEhJ6
niPxt9Ao6eG/7lV/NA9kvO58w6suGhdJYInMd7JRn/p/1Pes/amm/+7E83RROcUU
JqEOIvg0tlHtsSJUqlvy76YoRrDPk4EHCcYGJYorUo9I9g/+0KWt7Ck6VxTlcLRJ
vxTrdGC+dUoT5nV2ZN2Z/f7QskDXsuFD6ZCAp/qmTBIVEs9PIE5Hw9y+9m5U3Q42
GEiL1OXFhTeNAienxr/S02J5iT7yekdtsjJv+st+ibbOnvzL/FaC+4+4/+Ajp+ob
AXm6nKueAa7nUtRwzewSbVKwXTpK0nZPih23KOeGIt770JZXyvkCrLq2jkT9NK6R
TVmV4VUEWkRJML9zz2m2u7w+g/7zN8jcbitQ5BlX0r2tH9hSAD323xam0Pp65/JQ
5BR1QH292+qlERa96D0Hqe/buJu9lYFVCOQpDk+8oy7ASS4wJReeb18UIDoi2sWa
yA7rdvekF1rqRQeUtTADmWIkIJoEnPdaAQ3Kyu4ZpwUD8hseApiVpK5pIEPGhwes
SmcDi16zVFM1UprPibvGZQFVbCwtV+T/iaYwXdwBr018cBNlKtlxal6D3dtrvkKv
8lto0f0J2Exu32nwB4Nv1EhWAZ7NDJMAebW6YRiQojJH/WYMjcwHqpLVFP7qJIHH
GYjv5f7QGzXvA4obPPPl2CHIiJFr392EMw4uZfvies59xvFlmIRDnbgdX/yJA3YG
xdjSkFySeplfzkqKeExh60xtd96/UcDENRDHqfq/Ot4MkX8/JQXTjLDz+Y55yM7x
IeETeGgqhvr7MkGFgl4aRbVBH0V93NU7BkkQsoIijyVkn9ypLeSLFzJs/EPzf4FZ
1zfpQWSvVtsC4hcbjbUzViRziJK5MB0t72xSFnUFYSr4CBChlmmq6KTyH+gBq1ws
5nvOmiOLtgsY4npSumk3lIUvGkVlQpxco+cAMOZzny58HWPzXoWoLLS7C6AqoxUB
3/C77GeXMD+VonjvNYO4oA==
`pragma protect end_protected
